magic
tech sky130A
magscale 1 2
timestamp 1698067942
<< pwell >>
rect -246 -1179 246 1179
<< nmos >>
rect -50 -1031 50 969
<< ndiff >>
rect -108 957 -50 969
rect -108 -1019 -96 957
rect -62 -1019 -50 957
rect -108 -1031 -50 -1019
rect 50 957 108 969
rect 50 -1019 62 957
rect 96 -1019 108 957
rect 50 -1031 108 -1019
<< ndiffc >>
rect -96 -1019 -62 957
rect 62 -1019 96 957
<< psubdiff >>
rect -210 1109 210 1143
rect -210 -1109 -176 1109
rect 176 -1109 210 1109
rect -210 -1143 -114 -1109
rect 114 -1143 210 -1109
<< psubdiffcont >>
rect -114 -1143 114 -1109
<< poly >>
rect -50 1041 50 1057
rect -50 1007 -34 1041
rect 34 1007 50 1041
rect -50 969 50 1007
rect -50 -1057 50 -1031
<< polycont >>
rect -34 1007 34 1041
<< locali >>
rect -210 1109 210 1143
rect -210 -1109 -176 1109
rect -50 1007 -34 1041
rect 34 1007 50 1041
rect -96 957 -62 973
rect -96 -1035 -62 -1019
rect 62 957 96 973
rect 62 -1035 96 -1019
rect 176 -1109 210 1109
rect -210 -1143 -114 -1109
rect 114 -1143 210 -1109
<< properties >>
string FIXED_BBOX -193 -1126 193 1126
<< end >>
