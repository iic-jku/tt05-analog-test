magic
tech sky130A
magscale 1 2
timestamp 1698137664
<< locali >>
rect 4546 21109 4616 21115
rect 4546 21051 4551 21109
rect 4609 21051 4616 21109
rect 4546 20745 4616 21051
rect 5086 21109 5156 21113
rect 5086 21051 5091 21109
rect 5149 21051 5156 21109
rect 5086 20745 5156 21051
rect 5626 21109 5696 21111
rect 5626 21051 5631 21109
rect 5689 21051 5696 21109
rect 5626 20745 5696 21051
rect 6206 21109 6276 21111
rect 6206 21051 6211 21109
rect 6269 21051 6276 21109
rect 6206 20745 6276 21051
rect 6746 21109 6816 21111
rect 6746 21051 6751 21109
rect 6809 21051 6816 21109
rect 6746 20745 6816 21051
rect 7326 21109 7396 21111
rect 7326 21051 7327 21109
rect 7385 21051 7396 21109
rect 7326 20745 7396 21051
rect 7866 21109 7936 21113
rect 7866 21051 7871 21109
rect 7929 21051 7936 21109
rect 7866 20745 7936 21051
rect 8426 21109 8496 21111
rect 8426 21051 8431 21109
rect 8489 21051 8496 21109
rect 8426 20745 8496 21051
rect 8986 21109 9056 21113
rect 8986 21051 8991 21109
rect 9049 21051 9056 21109
rect 8986 20745 9056 21051
rect 9546 21109 9616 21115
rect 9546 21051 9551 21109
rect 9609 21051 9616 21109
rect 9546 20745 9616 21051
rect 10126 21109 10196 21115
rect 10126 21051 10131 21109
rect 10189 21051 10196 21109
rect 10126 20745 10196 21051
rect 10666 21109 10736 21113
rect 10666 21051 10671 21109
rect 10729 21051 10736 21109
rect 10666 20745 10736 21051
rect 11186 21109 11256 21115
rect 11186 21051 11191 21109
rect 11249 21051 11256 21109
rect 11186 20745 11256 21051
rect 11746 21109 11816 21113
rect 11746 21051 11751 21109
rect 11809 21051 11816 21109
rect 11746 20745 11816 21051
rect 12306 21109 12376 21115
rect 12306 21051 12311 21109
rect 12369 21051 12376 21109
rect 12306 20745 12376 21051
rect 12866 21109 12936 21115
rect 12866 21051 12871 21109
rect 12929 21051 12936 21109
rect 12866 20745 12936 21051
rect 13406 21109 13476 21115
rect 13406 21051 13411 21109
rect 13469 21051 13476 21109
rect 13406 20745 13476 21051
rect 13966 21109 14036 21111
rect 13966 21051 13971 21109
rect 14029 21051 14036 21109
rect 13966 20745 14036 21051
rect 14546 21109 14616 21113
rect 14546 21051 14551 21109
rect 14609 21051 14616 21109
rect 14546 20745 14616 21051
rect 15066 21109 15136 21115
rect 15066 21051 15071 21109
rect 15129 21051 15136 21109
rect 15066 20745 15136 21051
rect 15626 21109 15696 21117
rect 15626 21051 15631 21109
rect 15689 21051 15696 21109
rect 15626 20745 15696 21051
rect 16166 21109 16236 21113
rect 16166 21051 16171 21109
rect 16229 21051 16236 21109
rect 16166 20745 16236 21051
rect 16706 21109 16776 21119
rect 16706 21051 16711 21109
rect 16769 21051 16776 21109
rect 16706 20745 16776 21051
rect 17266 21109 17336 21113
rect 17266 21051 17271 21109
rect 17329 21051 17336 21109
rect 17266 20745 17336 21051
rect 14724 14534 15194 14536
rect 14260 14466 15194 14534
rect 14260 14464 14818 14466
rect 14256 12636 15530 12706
<< viali >>
rect 4551 21731 4609 21789
rect 5096 21736 5144 21784
rect 5636 21736 5684 21784
rect 6216 21736 6264 21784
rect 6756 21736 6804 21784
rect 7336 21736 7384 21784
rect 7876 21736 7924 21784
rect 8436 21736 8484 21784
rect 8996 21736 9044 21784
rect 9556 21736 9604 21784
rect 10136 21736 10184 21784
rect 10676 21736 10724 21784
rect 11196 21736 11244 21784
rect 11756 21736 11804 21784
rect 12316 21736 12364 21784
rect 12876 21736 12924 21784
rect 13416 21736 13464 21784
rect 13976 21736 14024 21784
rect 14556 21736 14604 21784
rect 15076 21736 15124 21784
rect 15636 21736 15684 21784
rect 16176 21736 16224 21784
rect 16716 21736 16764 21784
rect 17276 21736 17324 21784
rect 4551 21051 4609 21109
rect 5091 21051 5149 21109
rect 5631 21051 5689 21109
rect 6211 21051 6269 21109
rect 6751 21051 6809 21109
rect 7327 21051 7385 21109
rect 7871 21051 7929 21109
rect 8431 21051 8489 21109
rect 8991 21051 9049 21109
rect 9551 21051 9609 21109
rect 10131 21051 10189 21109
rect 10671 21051 10729 21109
rect 11191 21051 11249 21109
rect 11751 21051 11809 21109
rect 12311 21051 12369 21109
rect 12871 21051 12929 21109
rect 13411 21051 13469 21109
rect 13971 21051 14029 21109
rect 14551 21051 14609 21109
rect 15071 21051 15129 21109
rect 15631 21051 15689 21109
rect 16171 21051 16229 21109
rect 16711 21051 16769 21109
rect 17271 21051 17329 21109
rect 18955 16543 18989 16577
rect 19447 16543 19481 16577
rect 19939 16533 19973 16569
rect 18875 15479 18909 15513
rect 19367 15479 19401 15513
rect 19859 15479 19893 15513
rect 12975 15035 13009 15069
rect 13467 15035 13501 15069
rect 13959 15035 13993 15069
rect 12895 14471 12929 14505
rect 13387 14471 13421 14505
rect 13879 14479 13913 14513
rect 19033 14491 19067 14525
rect 19525 14491 19559 14525
rect 20017 14491 20051 14525
rect 18841 14383 18875 14417
rect 19333 14383 19367 14417
rect 19825 14383 19859 14417
rect 14587 14317 14621 14351
rect 15299 14317 15333 14351
rect 14587 14151 14621 14185
rect 15299 14151 15333 14185
rect 19207 14167 19241 14201
rect 19875 14165 19909 14199
rect 18911 14087 18945 14121
rect 19471 14087 19505 14121
rect 19681 14085 19715 14119
rect 20031 14085 20065 14119
rect 13053 13983 13087 14017
rect 13545 13983 13579 14017
rect 14037 13993 14071 14027
rect 14587 13985 14621 14019
rect 15299 13985 15333 14019
rect 19019 14007 19053 14041
rect 19789 14007 19823 14041
rect 12975 13875 13009 13909
rect 13467 13875 13501 13909
rect 13959 13887 13993 13921
rect 14587 13819 14621 13853
rect 15299 13819 15333 13853
rect 12975 13771 13009 13805
rect 13467 13771 13501 13805
rect 13959 13779 13993 13813
rect 16879 13763 16913 13797
rect 17687 13765 17721 13799
rect 12897 13663 12931 13697
rect 13389 13663 13423 13697
rect 13881 13673 13915 13707
rect 14587 13653 14621 13687
rect 15299 13653 15333 13687
rect 15835 13685 15869 13719
rect 16987 13685 17021 13719
rect 17091 13685 17125 13719
rect 18243 13685 18277 13719
rect 16391 13605 16425 13639
rect 17199 13607 17233 13641
rect 14257 13569 14291 13603
rect 14587 13487 14621 13521
rect 15299 13487 15333 13521
rect 19107 13419 19141 13453
rect 19877 13417 19911 13451
rect 14587 13321 14621 13355
rect 15299 13321 15333 13355
rect 18865 13339 18899 13373
rect 19215 13339 19249 13373
rect 19425 13339 19459 13373
rect 19985 13339 20019 13373
rect 16891 13271 16925 13305
rect 17699 13273 17733 13307
rect 19021 13259 19055 13293
rect 19689 13259 19723 13293
rect 13055 13175 13089 13209
rect 13547 13175 13581 13209
rect 14039 13187 14073 13221
rect 15839 13193 15873 13227
rect 16999 13193 17033 13227
rect 17103 13193 17137 13227
rect 18263 13193 18297 13227
rect 14587 13155 14621 13189
rect 15299 13155 15333 13189
rect 16403 13113 16437 13147
rect 17211 13115 17245 13149
rect 19071 13041 19105 13075
rect 19563 13041 19597 13075
rect 20055 13041 20089 13075
rect 14587 12989 14621 13023
rect 15299 12989 15333 13023
rect 18879 12935 18913 12969
rect 19371 12933 19405 12967
rect 19863 12933 19897 12967
rect 14587 12823 14621 12857
rect 15299 12823 15333 12857
rect 16891 12779 16925 12813
rect 17699 12781 17733 12815
rect 12975 12611 13009 12645
rect 13467 12611 13501 12645
rect 13959 12631 13993 12665
rect 15839 12701 15873 12735
rect 16999 12701 17033 12735
rect 17103 12701 17137 12735
rect 18263 12701 18297 12735
rect 16403 12621 16437 12655
rect 17211 12623 17245 12657
rect 13937 12031 13971 12065
rect 14745 12035 14779 12069
rect 16917 12033 16951 12067
rect 17723 12035 17757 12069
rect 12885 11955 12919 11989
rect 14045 11955 14079 11989
rect 14149 11955 14183 11989
rect 15309 11955 15343 11989
rect 15873 11955 15907 11989
rect 17023 11955 17057 11989
rect 17129 11955 17163 11989
rect 18279 11955 18313 11989
rect 19037 11947 19071 11981
rect 19529 11945 19563 11979
rect 20021 11945 20055 11979
rect 13449 11875 13483 11909
rect 14257 11875 14291 11909
rect 16429 11875 16463 11909
rect 17237 11877 17271 11911
rect 13937 11539 13971 11573
rect 14745 11543 14779 11577
rect 16927 11541 16961 11575
rect 17735 11543 17769 11577
rect 12885 11463 12919 11497
rect 14045 11463 14079 11497
rect 14149 11463 14183 11497
rect 15309 11463 15343 11497
rect 15875 11463 15909 11497
rect 17035 11463 17069 11497
rect 17139 11463 17173 11497
rect 18299 11463 18333 11497
rect 13449 11383 13483 11417
rect 14257 11383 14291 11417
rect 16439 11383 16473 11417
rect 17247 11385 17281 11419
rect 13947 11047 13981 11081
rect 14755 11051 14789 11085
rect 16927 11049 16961 11083
rect 17735 11051 17769 11085
rect 12905 10971 12939 11005
rect 14055 10971 14089 11005
rect 14161 10971 14195 11005
rect 15311 10971 15345 11005
rect 15875 10971 15909 11005
rect 17035 10971 17069 11005
rect 17139 10971 17173 11005
rect 18299 10971 18333 11005
rect 13461 10891 13495 10925
rect 14267 10891 14301 10925
rect 16439 10891 16473 10925
rect 17247 10893 17281 10927
rect 18957 10891 18991 10925
rect 19449 10881 19483 10915
rect 19941 10881 19975 10915
rect 13229 10315 13263 10349
rect 13721 10315 13755 10349
rect 14213 10303 14247 10337
rect 13149 9251 13183 9285
rect 13641 9251 13675 9285
rect 14133 9247 14167 9281
rect 19068 8916 19334 9470
rect 18157 8793 18191 8827
rect 17063 8713 17097 8747
rect 19213 8713 19247 8747
rect 17171 8633 17205 8667
rect 18147 8301 18181 8335
rect 13307 8263 13341 8297
rect 13799 8263 13833 8297
rect 14291 8261 14325 8295
rect 17051 8221 17085 8255
rect 19211 8221 19245 8255
rect 13115 8155 13149 8189
rect 13607 8155 13641 8189
rect 14099 8155 14133 8189
rect 17159 8141 17193 8175
rect 13481 7935 13515 7969
rect 14149 7935 14183 7969
rect 13185 7855 13219 7889
rect 13745 7855 13779 7889
rect 13955 7855 13989 7889
rect 14305 7855 14339 7889
rect 13293 7779 13327 7813
rect 14061 7777 14095 7811
rect 18147 7809 18181 7843
rect 17051 7729 17085 7763
rect 19211 7729 19245 7763
rect 17159 7649 17193 7683
rect 14973 7301 15007 7335
rect 13879 7221 13913 7255
rect 16029 7221 16063 7255
rect 13987 7143 14021 7177
rect 19209 7061 19243 7095
rect 17157 6933 17191 6967
rect 19317 6933 19351 6967
rect 14963 6809 14997 6843
rect 18221 6801 18255 6835
rect 13867 6729 13901 6763
rect 16027 6729 16061 6763
rect 13975 6651 14009 6685
rect 16581 6481 16615 6515
rect 18173 6481 18207 6515
rect 17143 6365 17177 6399
rect 14963 6317 14997 6351
rect 19201 6329 19235 6363
rect 13867 6237 13901 6271
rect 16027 6237 16061 6271
rect 18173 6221 18207 6255
rect 13975 6159 14009 6193
rect 19209 6001 19243 6035
rect 17157 5773 17191 5807
rect 19317 5773 19351 5807
rect 13277 5685 13311 5719
rect 14437 5685 14471 5719
rect 13149 5577 13183 5611
rect 13881 5569 13915 5603
rect 14209 5577 14243 5611
rect 15131 5569 15165 5603
rect 15489 5571 15523 5605
rect 18221 5541 18255 5575
rect 16351 5425 16385 5459
rect 18173 5221 18207 5255
rect 17143 5115 17177 5149
rect 19201 5077 19235 5111
rect 17109 4971 17143 5005
rect 18173 4865 18207 4899
rect 17145 4757 17179 4791
rect 19203 4721 19237 4755
rect 13407 4589 13441 4623
rect 14667 4589 14701 4623
rect 18173 4615 18207 4649
rect 13729 4541 13763 4575
rect 13989 4541 14023 4575
rect 14989 4541 15023 4575
rect 15345 4541 15379 4575
rect 15595 4541 15629 4575
rect 16809 4439 16843 4473
rect 16581 4333 16615 4367
rect 18973 4225 19007 4259
rect 18745 4119 18779 4153
rect 17381 3943 17415 3977
rect 16351 3837 16385 3871
rect 18409 3801 18443 3835
rect 17381 3693 17415 3727
rect 18445 3587 18479 3621
rect 13277 3525 13311 3559
rect 13843 3511 13877 3545
rect 14437 3525 14471 3559
rect 15095 3511 15129 3545
rect 15451 3513 15485 3547
rect 15239 3477 15273 3511
rect 16353 3481 16387 3515
rect 18411 3443 18445 3477
rect 17381 3337 17415 3371
rect 15771 3177 15805 3211
rect 19203 3133 19237 3167
rect 17333 3017 17367 3051
rect 13727 2949 13761 2983
rect 15877 2949 15911 2983
rect 16237 2785 16271 2819
rect 18397 2785 18431 2819
rect 14783 2719 14817 2753
rect 16345 2557 16379 2591
rect 14719 2387 14753 2421
rect 13625 2307 13659 2341
rect 15775 2307 15809 2341
rect 17381 2337 17415 2371
rect 13733 2229 13767 2263
rect 16353 2229 16387 2263
rect 18411 2193 18445 2227
rect 17381 2077 17415 2111
rect 18973 2077 19007 2111
rect 14709 1895 14743 1929
rect 13613 1815 13647 1849
rect 15773 1815 15807 1849
rect 13721 1737 13755 1771
rect 17333 1757 17367 1791
rect 16237 1625 16271 1659
rect 18397 1625 18431 1659
rect 16345 1497 16379 1531
rect 14709 1403 14743 1437
rect 13613 1323 13647 1357
rect 15773 1323 15807 1357
rect 13721 1245 13755 1279
<< metal1 >>
rect 5060 22251 5180 22280
rect 4539 22145 4545 22215
rect 4615 22145 4621 22215
rect 5060 22191 5090 22251
rect 5150 22191 5180 22251
rect 5060 22160 5180 22191
rect 5600 22250 5720 22280
rect 5600 22190 5630 22250
rect 5690 22190 5720 22250
rect 5600 22160 5720 22190
rect 6180 22250 6300 22280
rect 6180 22190 6210 22250
rect 6270 22190 6300 22250
rect 6180 22160 6300 22190
rect 6720 22250 6840 22280
rect 6720 22190 6750 22250
rect 6810 22190 6840 22250
rect 6720 22160 6840 22190
rect 7300 22250 7420 22280
rect 7300 22190 7330 22250
rect 7390 22190 7420 22250
rect 7300 22160 7420 22190
rect 7840 22250 7960 22280
rect 7840 22190 7870 22250
rect 7930 22190 7960 22250
rect 7840 22160 7960 22190
rect 8400 22250 8520 22280
rect 8400 22190 8430 22250
rect 8490 22190 8520 22250
rect 8400 22160 8520 22190
rect 8960 22250 9080 22280
rect 8960 22190 8990 22250
rect 9050 22190 9080 22250
rect 8960 22160 9080 22190
rect 9520 22250 9640 22280
rect 9520 22190 9550 22250
rect 9610 22190 9640 22250
rect 9520 22160 9640 22190
rect 10100 22250 10220 22280
rect 10100 22190 10130 22250
rect 10190 22190 10220 22250
rect 10100 22160 10220 22190
rect 10640 22250 10760 22280
rect 10640 22190 10670 22250
rect 10730 22190 10760 22250
rect 10640 22160 10760 22190
rect 11160 22250 11280 22280
rect 11160 22190 11190 22250
rect 11250 22190 11280 22250
rect 11160 22160 11280 22190
rect 11720 22250 11840 22280
rect 11720 22190 11750 22250
rect 11810 22190 11840 22250
rect 11720 22160 11840 22190
rect 12280 22250 12400 22280
rect 12280 22190 12310 22250
rect 12370 22190 12400 22250
rect 12280 22160 12400 22190
rect 12840 22250 12960 22280
rect 12840 22190 12870 22250
rect 12930 22190 12960 22250
rect 12840 22160 12960 22190
rect 13380 22250 13500 22280
rect 13380 22190 13410 22250
rect 13470 22190 13500 22250
rect 13380 22160 13500 22190
rect 13940 22250 14060 22280
rect 13940 22190 13970 22250
rect 14030 22190 14060 22250
rect 13940 22160 14060 22190
rect 14520 22250 14640 22280
rect 14520 22190 14550 22250
rect 14610 22190 14640 22250
rect 14520 22160 14640 22190
rect 15040 22250 15160 22280
rect 15040 22190 15070 22250
rect 15130 22190 15160 22250
rect 15040 22160 15160 22190
rect 15600 22250 15720 22280
rect 15600 22190 15630 22250
rect 15690 22190 15720 22250
rect 15600 22160 15720 22190
rect 16140 22250 16260 22280
rect 16140 22190 16170 22250
rect 16230 22190 16260 22250
rect 16140 22160 16260 22190
rect 16680 22250 16800 22280
rect 16680 22190 16710 22250
rect 16770 22190 16800 22250
rect 16680 22160 16800 22190
rect 17240 22250 17360 22280
rect 17240 22190 17270 22250
rect 17330 22190 17360 22250
rect 17240 22160 17360 22190
rect 4545 21789 4615 22145
rect 4545 21731 4551 21789
rect 4609 21731 4615 21789
rect 4545 21719 4615 21731
rect 5090 21784 5150 22160
rect 5090 21736 5096 21784
rect 5144 21736 5150 21784
rect 5090 21724 5150 21736
rect 5630 21784 5690 22160
rect 5630 21736 5636 21784
rect 5684 21736 5690 21784
rect 5630 21724 5690 21736
rect 6210 21784 6270 22160
rect 6210 21736 6216 21784
rect 6264 21736 6270 21784
rect 6210 21724 6270 21736
rect 6750 21784 6810 22160
rect 6750 21736 6756 21784
rect 6804 21736 6810 21784
rect 6750 21724 6810 21736
rect 7330 21784 7390 22160
rect 7330 21736 7336 21784
rect 7384 21736 7390 21784
rect 7330 21724 7390 21736
rect 7870 21784 7930 22160
rect 7870 21736 7876 21784
rect 7924 21736 7930 21784
rect 7870 21724 7930 21736
rect 8430 21784 8490 22160
rect 8430 21736 8436 21784
rect 8484 21736 8490 21784
rect 8430 21724 8490 21736
rect 8990 21784 9050 22160
rect 8990 21736 8996 21784
rect 9044 21736 9050 21784
rect 8990 21724 9050 21736
rect 9550 21784 9610 22160
rect 9550 21736 9556 21784
rect 9604 21736 9610 21784
rect 9550 21724 9610 21736
rect 10130 21784 10190 22160
rect 10130 21736 10136 21784
rect 10184 21736 10190 21784
rect 10130 21724 10190 21736
rect 10670 21784 10730 22160
rect 10670 21736 10676 21784
rect 10724 21736 10730 21784
rect 10670 21724 10730 21736
rect 11190 21784 11250 22160
rect 11190 21736 11196 21784
rect 11244 21736 11250 21784
rect 11190 21724 11250 21736
rect 11750 21784 11810 22160
rect 11750 21736 11756 21784
rect 11804 21736 11810 21784
rect 11750 21724 11810 21736
rect 12310 21784 12370 22160
rect 12310 21736 12316 21784
rect 12364 21736 12370 21784
rect 12310 21724 12370 21736
rect 12870 21784 12930 22160
rect 12870 21736 12876 21784
rect 12924 21736 12930 21784
rect 12870 21724 12930 21736
rect 13410 21784 13470 22160
rect 13410 21736 13416 21784
rect 13464 21736 13470 21784
rect 13410 21724 13470 21736
rect 13970 21784 14030 22160
rect 13970 21736 13976 21784
rect 14024 21736 14030 21784
rect 13970 21724 14030 21736
rect 14550 21784 14610 22160
rect 14550 21736 14556 21784
rect 14604 21736 14610 21784
rect 14550 21724 14610 21736
rect 15070 21784 15130 22160
rect 15070 21736 15076 21784
rect 15124 21736 15130 21784
rect 15070 21724 15130 21736
rect 15630 21784 15690 22160
rect 15630 21736 15636 21784
rect 15684 21736 15690 21784
rect 15630 21724 15690 21736
rect 16170 21784 16230 22160
rect 16170 21736 16176 21784
rect 16224 21736 16230 21784
rect 16170 21724 16230 21736
rect 16710 21784 16770 22160
rect 16710 21736 16716 21784
rect 16764 21736 16770 21784
rect 16710 21724 16770 21736
rect 17270 21784 17330 22160
rect 17270 21736 17276 21784
rect 17324 21736 17330 21784
rect 17270 21724 17330 21736
rect 18952 21115 18958 21120
rect 4525 21109 18958 21115
rect 4525 21051 4551 21109
rect 4609 21051 5091 21109
rect 5149 21051 5631 21109
rect 5689 21051 6211 21109
rect 6269 21051 6751 21109
rect 6809 21051 7327 21109
rect 7385 21051 7871 21109
rect 7929 21051 8431 21109
rect 8489 21051 8991 21109
rect 9049 21051 9551 21109
rect 9609 21051 10131 21109
rect 10189 21051 10671 21109
rect 10729 21051 11191 21109
rect 11249 21051 11751 21109
rect 11809 21051 12311 21109
rect 12369 21051 12871 21109
rect 12929 21051 13411 21109
rect 13469 21051 13971 21109
rect 14029 21051 14551 21109
rect 14609 21051 15071 21109
rect 15129 21051 15631 21109
rect 15689 21051 16171 21109
rect 16229 21051 16711 21109
rect 16769 21051 17271 21109
rect 17329 21051 18958 21109
rect 4525 21045 18958 21051
rect 18952 21035 18958 21045
rect 19043 21115 19049 21120
rect 19043 21045 19051 21115
rect 19043 21035 19049 21045
rect 19838 16650 20070 16672
rect 18943 16577 19001 16589
rect 18943 16543 18955 16577
rect 18989 16574 19001 16577
rect 19190 16574 19196 16586
rect 18989 16546 19196 16574
rect 18989 16543 19001 16546
rect 18943 16531 19001 16543
rect 19190 16534 19196 16546
rect 19248 16574 19254 16586
rect 19435 16577 19493 16589
rect 19435 16574 19447 16577
rect 19248 16546 19447 16574
rect 19248 16534 19254 16546
rect 19435 16543 19447 16546
rect 19481 16543 19493 16577
rect 19435 16531 19493 16543
rect 19838 16450 19860 16650
rect 20050 16450 20070 16650
rect 19838 16430 20070 16450
rect 18863 15513 18921 15525
rect 18863 15479 18875 15513
rect 18909 15510 18921 15513
rect 19349 15522 19423 15533
rect 19349 15510 19360 15522
rect 18909 15482 19360 15510
rect 18909 15479 18921 15482
rect 18863 15467 18921 15479
rect 19349 15470 19360 15482
rect 19412 15510 19423 15522
rect 19847 15513 19905 15525
rect 19847 15510 19859 15513
rect 19412 15482 19859 15510
rect 19412 15470 19423 15482
rect 19349 15459 19423 15470
rect 19847 15479 19859 15482
rect 19893 15479 19905 15513
rect 19847 15467 19905 15479
rect 12963 15069 13021 15081
rect 12963 15035 12975 15069
rect 13009 15066 13021 15069
rect 13455 15069 13513 15081
rect 13455 15066 13467 15069
rect 13009 15038 13467 15066
rect 13009 15035 13021 15038
rect 12963 15023 13021 15035
rect 13455 15035 13467 15038
rect 13501 15066 13513 15069
rect 13947 15069 14005 15081
rect 13947 15066 13959 15069
rect 13501 15038 13959 15066
rect 13501 15035 13513 15038
rect 13455 15023 13513 15035
rect 13947 15035 13959 15038
rect 13993 15066 14005 15069
rect 13993 15035 14006 15066
rect 13947 15023 14006 15035
rect 12883 14505 12941 14517
rect 12883 14471 12895 14505
rect 12929 14502 12941 14505
rect 13375 14510 13433 14517
rect 13867 14513 13925 14525
rect 13867 14510 13879 14513
rect 13375 14505 13879 14510
rect 13375 14502 13387 14505
rect 12929 14474 13387 14502
rect 12929 14471 12941 14474
rect 12883 14459 12941 14471
rect 13375 14471 13387 14474
rect 13421 14482 13879 14505
rect 13421 14471 13433 14482
rect 13375 14459 13433 14471
rect 13867 14479 13879 14482
rect 13913 14479 13925 14513
rect 13867 14467 13925 14479
rect 13882 14371 13910 14467
rect 13875 14360 13949 14371
rect 13875 14308 13886 14360
rect 13938 14308 13949 14360
rect 13875 14297 13949 14308
rect 13978 14149 14006 15023
rect 19021 14525 19079 14537
rect 19021 14522 19033 14525
rect 15222 14494 19033 14522
rect 14035 14360 14109 14371
rect 14035 14308 14046 14360
rect 14098 14348 14109 14360
rect 14575 14351 14633 14363
rect 14575 14348 14587 14351
rect 14098 14320 14587 14348
rect 14098 14308 14109 14320
rect 14035 14297 14109 14308
rect 14575 14317 14587 14320
rect 14621 14317 14633 14351
rect 14575 14305 14633 14317
rect 15222 14276 15250 14494
rect 19021 14491 19033 14494
rect 19067 14522 19079 14525
rect 19505 14534 19579 14545
rect 19505 14522 19516 14534
rect 19067 14494 19516 14522
rect 19067 14491 19079 14494
rect 19021 14479 19079 14491
rect 19505 14482 19516 14494
rect 19568 14482 19579 14534
rect 19505 14471 19579 14482
rect 18829 14417 18887 14429
rect 18829 14383 18841 14417
rect 18875 14414 18887 14417
rect 19322 14417 19382 14430
rect 19823 14429 19897 14437
rect 19322 14414 19333 14417
rect 18875 14386 19333 14414
rect 18875 14383 18887 14386
rect 18829 14371 18887 14383
rect 19322 14383 19333 14386
rect 19367 14383 19382 14417
rect 15287 14351 15345 14363
rect 15287 14317 15299 14351
rect 15333 14317 15345 14351
rect 15287 14305 15345 14317
rect 14590 14248 15250 14276
rect 14590 14197 14618 14248
rect 15302 14197 15330 14305
rect 14575 14185 14633 14197
rect 14575 14151 14587 14185
rect 14621 14151 14633 14185
rect 13955 14138 14029 14149
rect 14575 14139 14633 14151
rect 15287 14185 15345 14197
rect 15287 14151 15299 14185
rect 15333 14151 15345 14185
rect 15287 14139 15345 14151
rect 13955 14086 13966 14138
rect 14018 14086 14029 14138
rect 13955 14075 14029 14086
rect 13041 14017 13099 14029
rect 13041 14014 13053 14017
rect 12978 13986 13053 14014
rect 12978 13921 13006 13986
rect 13041 13983 13053 13986
rect 13087 13983 13099 14017
rect 13041 13971 13099 13983
rect 13533 14017 13591 14029
rect 14025 14027 14083 14039
rect 14590 14031 14618 14139
rect 18844 14134 18872 14371
rect 19322 14370 19382 14383
rect 19813 14426 19897 14429
rect 19813 14417 19834 14426
rect 19813 14383 19825 14417
rect 19813 14374 19834 14383
rect 19886 14374 19897 14426
rect 19813 14371 19897 14374
rect 19823 14363 19897 14371
rect 18963 14346 19037 14357
rect 18963 14294 18974 14346
rect 19026 14334 19037 14346
rect 19026 14306 19122 14334
rect 19026 14294 19037 14306
rect 18963 14283 19037 14294
rect 18844 14121 18958 14134
rect 18844 14087 18911 14121
rect 18945 14118 18958 14121
rect 18945 14090 19050 14118
rect 18945 14087 18958 14090
rect 18844 14074 18958 14087
rect 19022 14053 19050 14090
rect 19007 14041 19065 14053
rect 14025 14024 14037 14027
rect 13533 13983 13545 14017
rect 13579 13983 13591 14017
rect 13533 13971 13591 13983
rect 13962 13996 14037 14024
rect 12963 13909 13021 13921
rect 12963 13875 12975 13909
rect 13009 13875 13021 13909
rect 12963 13863 13021 13875
rect 13455 13909 13513 13921
rect 13455 13875 13467 13909
rect 13501 13906 13513 13909
rect 13548 13906 13576 13971
rect 13962 13933 13990 13996
rect 14025 13993 14037 13996
rect 14071 13993 14083 14027
rect 14025 13981 14083 13993
rect 14575 14019 14633 14031
rect 14575 13985 14587 14019
rect 14621 13985 14633 14019
rect 14575 13973 14633 13985
rect 15287 14019 15345 14031
rect 15287 13985 15299 14019
rect 15333 13985 15345 14019
rect 19007 14007 19019 14041
rect 19053 14007 19065 14041
rect 19094 14038 19122 14306
rect 19942 14268 19970 16430
rect 19999 14534 20073 14545
rect 19999 14482 20010 14534
rect 20062 14482 20073 14534
rect 19999 14471 20073 14482
rect 19942 14240 19978 14268
rect 19188 14208 19258 14222
rect 19188 14156 19196 14208
rect 19248 14156 19258 14208
rect 19823 14211 19897 14219
rect 19823 14208 19921 14211
rect 19188 14142 19258 14156
rect 19458 14160 19786 14188
rect 19458 14121 19518 14160
rect 19458 14087 19471 14121
rect 19505 14087 19518 14121
rect 19458 14074 19518 14087
rect 19669 14119 19727 14131
rect 19669 14085 19681 14119
rect 19715 14085 19727 14119
rect 19758 14116 19786 14160
rect 19823 14156 19834 14208
rect 19886 14199 19921 14208
rect 19909 14165 19921 14199
rect 19886 14156 19921 14165
rect 19823 14153 19921 14156
rect 19823 14145 19897 14153
rect 19950 14116 19978 14240
rect 20019 14119 20077 14131
rect 20019 14116 20031 14119
rect 19758 14088 20031 14116
rect 19669 14073 19727 14085
rect 20019 14085 20031 14088
rect 20065 14085 20077 14119
rect 20019 14073 20077 14085
rect 19684 14038 19712 14073
rect 19769 14048 19843 14059
rect 19769 14038 19780 14048
rect 19094 14010 19780 14038
rect 19007 13995 19065 14007
rect 15287 13973 15345 13985
rect 13501 13878 13576 13906
rect 13947 13921 14005 13933
rect 13947 13887 13959 13921
rect 13993 13887 14005 13921
rect 13501 13875 13513 13878
rect 13947 13875 14005 13887
rect 13455 13863 13513 13875
rect 12978 13817 13006 13863
rect 13470 13817 13498 13863
rect 13962 13825 13990 13875
rect 15302 13865 15330 13973
rect 18146 13947 18382 13960
rect 14575 13853 14633 13865
rect 12963 13805 13021 13817
rect 12963 13802 12975 13805
rect 12900 13774 12975 13802
rect 12900 13709 12928 13774
rect 12963 13771 12975 13774
rect 13009 13771 13021 13805
rect 12963 13759 13021 13771
rect 13455 13805 13513 13817
rect 13947 13813 14005 13825
rect 13947 13810 13959 13813
rect 13455 13771 13467 13805
rect 13501 13771 13513 13805
rect 13455 13759 13513 13771
rect 13884 13782 13959 13810
rect 12885 13697 12943 13709
rect 12885 13663 12897 13697
rect 12931 13694 12943 13697
rect 13377 13697 13435 13709
rect 13377 13694 13389 13697
rect 12931 13674 13389 13694
rect 13423 13694 13435 13697
rect 13470 13694 13498 13759
rect 13884 13719 13912 13782
rect 13947 13779 13959 13782
rect 13993 13779 14005 13813
rect 14575 13819 14587 13853
rect 14621 13819 14633 13853
rect 14575 13807 14633 13819
rect 15287 13853 15345 13865
rect 15287 13819 15299 13853
rect 15333 13819 15345 13853
rect 15287 13807 15345 13819
rect 13947 13767 14005 13779
rect 14590 13764 14618 13807
rect 13955 13728 14029 13739
rect 14590 13736 15250 13764
rect 13423 13674 13498 13694
rect 12885 13651 12914 13663
rect 12904 13444 12914 13651
rect 13478 13444 13498 13674
rect 13869 13707 13927 13719
rect 13869 13673 13881 13707
rect 13915 13673 13927 13707
rect 13869 13661 13927 13673
rect 13955 13676 13966 13728
rect 14018 13676 14029 13728
rect 13955 13665 14029 13676
rect 14575 13687 14633 13699
rect 13884 13623 13912 13661
rect 13859 13612 13933 13623
rect 13859 13560 13870 13612
rect 13922 13560 13933 13612
rect 13859 13549 13933 13560
rect 13470 13323 13498 13444
rect 13447 13312 13521 13323
rect 13447 13260 13458 13312
rect 13510 13260 13521 13312
rect 13447 13249 13521 13260
rect 13043 13209 13101 13221
rect 13043 13175 13055 13209
rect 13089 13206 13101 13209
rect 13535 13218 13593 13221
rect 13962 13218 13990 13665
rect 14575 13653 14587 13687
rect 14621 13653 14633 13687
rect 14575 13641 14633 13653
rect 14019 13612 14093 13623
rect 14019 13560 14030 13612
rect 14082 13600 14093 13612
rect 14245 13603 14303 13615
rect 14245 13600 14257 13603
rect 14082 13572 14257 13600
rect 14082 13560 14093 13572
rect 14019 13549 14093 13560
rect 14245 13569 14257 13572
rect 14291 13600 14303 13603
rect 14435 13612 14509 13623
rect 14435 13600 14446 13612
rect 14291 13572 14446 13600
rect 14291 13569 14303 13572
rect 14245 13557 14303 13569
rect 14435 13560 14446 13572
rect 14498 13560 14509 13612
rect 14435 13549 14509 13560
rect 14590 13533 14618 13641
rect 14575 13521 14633 13533
rect 14575 13487 14587 13521
rect 14621 13487 14633 13521
rect 14575 13475 14633 13487
rect 14575 13355 14633 13367
rect 14575 13321 14587 13355
rect 14621 13321 14633 13355
rect 15222 13352 15250 13736
rect 15302 13699 15330 13807
rect 16867 13797 16925 13809
rect 16867 13763 16879 13797
rect 16913 13763 16925 13797
rect 16867 13751 16925 13763
rect 17675 13799 17733 13811
rect 17675 13765 17687 13799
rect 17721 13765 17733 13799
rect 17675 13753 17733 13765
rect 15823 13719 15881 13731
rect 15287 13687 15345 13699
rect 15287 13653 15299 13687
rect 15333 13653 15345 13687
rect 15823 13685 15835 13719
rect 15869 13685 15881 13719
rect 16882 13716 16910 13751
rect 16974 13719 17034 13732
rect 16974 13716 16987 13719
rect 16882 13688 16987 13716
rect 15823 13673 15881 13685
rect 16920 13685 16987 13688
rect 17021 13716 17034 13719
rect 17079 13719 17137 13731
rect 17079 13716 17091 13719
rect 17021 13688 17091 13716
rect 17021 13685 17034 13688
rect 15287 13641 15345 13653
rect 15286 13530 15436 13542
rect 15286 13521 15372 13530
rect 15286 13487 15299 13521
rect 15333 13487 15372 13521
rect 15286 13478 15372 13487
rect 15424 13478 15436 13530
rect 15286 13466 15436 13478
rect 15278 13364 15354 13370
rect 15278 13352 15290 13364
rect 15222 13324 15290 13352
rect 14575 13309 14633 13321
rect 15278 13312 15290 13324
rect 15342 13312 15354 13364
rect 14027 13221 14085 13233
rect 14027 13218 14039 13221
rect 13535 13209 14039 13218
rect 13535 13206 13547 13209
rect 13089 13178 13547 13206
rect 13089 13175 13101 13178
rect 13043 13163 13101 13175
rect 13535 13175 13547 13178
rect 13581 13190 14039 13209
rect 13581 13175 13593 13190
rect 14027 13187 14039 13190
rect 14073 13187 14085 13221
rect 14590 13201 14618 13309
rect 15278 13308 15354 13312
rect 15842 13239 15870 13673
rect 16920 13672 17034 13685
rect 17079 13685 17091 13688
rect 17125 13716 17137 13719
rect 17125 13688 17230 13716
rect 17125 13685 17137 13688
rect 17079 13673 17137 13685
rect 16379 13639 16437 13651
rect 16379 13605 16391 13639
rect 16425 13605 16437 13639
rect 16379 13593 16437 13605
rect 16481 13612 16555 13623
rect 15899 13530 15973 13541
rect 15899 13478 15910 13530
rect 15962 13518 15973 13530
rect 16394 13518 16422 13593
rect 16481 13560 16492 13612
rect 16544 13600 16555 13612
rect 16920 13600 16948 13672
rect 17202 13653 17230 13688
rect 16544 13572 16948 13600
rect 17187 13641 17245 13653
rect 17187 13607 17199 13641
rect 17233 13607 17245 13641
rect 17187 13595 17245 13607
rect 16544 13560 16555 13572
rect 16481 13549 16555 13560
rect 15962 13490 16422 13518
rect 15962 13478 15973 13490
rect 15899 13467 15973 13478
rect 15827 13227 15885 13239
rect 14027 13175 14085 13187
rect 14575 13189 14633 13201
rect 13535 13163 13593 13175
rect 14575 13155 14587 13189
rect 14621 13155 14633 13189
rect 15287 13189 15345 13201
rect 15287 13186 15299 13189
rect 14575 13143 14633 13155
rect 15190 13158 15299 13186
rect 13927 13110 14001 13121
rect 13927 13058 13938 13110
rect 13990 13058 14001 13110
rect 13927 13047 14001 13058
rect 13950 12779 13978 13047
rect 14575 13023 14633 13035
rect 14575 12989 14587 13023
rect 14621 12989 14633 13023
rect 14575 12977 14633 12989
rect 14590 12869 14618 12977
rect 14575 12857 14633 12869
rect 14575 12823 14587 12857
rect 14621 12823 14633 12857
rect 14575 12811 14633 12823
rect 13927 12768 14001 12779
rect 12840 12645 13080 12730
rect 13927 12716 13938 12768
rect 13990 12716 14001 12768
rect 13927 12705 14001 12716
rect 13947 12665 14005 12677
rect 13947 12662 13959 12665
rect 13470 12657 13959 12662
rect 12840 12611 12975 12645
rect 13009 12642 13080 12645
rect 13455 12645 13959 12657
rect 13455 12642 13467 12645
rect 13009 12614 13467 12642
rect 13009 12611 13080 12614
rect 12840 12492 13080 12611
rect 13455 12611 13467 12614
rect 13501 12634 13959 12645
rect 13501 12611 13513 12634
rect 13947 12631 13959 12634
rect 13993 12631 14005 12665
rect 13947 12619 14005 12631
rect 13455 12599 13513 12611
rect 12816 12470 13154 12492
rect 12816 12230 12840 12470
rect 13080 12230 13154 12470
rect 12816 12194 13154 12230
rect 13447 12158 13521 12169
rect 13447 12106 13458 12158
rect 13510 12146 13521 12158
rect 13510 12118 13968 12146
rect 13510 12106 13521 12118
rect 13447 12095 13521 12106
rect 12873 11989 12931 12001
rect 12873 11955 12885 11989
rect 12919 11955 12931 11989
rect 12873 11943 12931 11955
rect 12888 11509 12916 11943
rect 13437 11909 13495 11921
rect 13437 11875 13449 11909
rect 13483 11875 13495 11909
rect 13437 11863 13495 11875
rect 12873 11497 12931 11509
rect 12873 11463 12885 11497
rect 12919 11494 12931 11497
rect 12919 11463 12936 11494
rect 12873 11451 12936 11463
rect 12908 11017 12936 11451
rect 13452 11429 13480 11863
rect 13437 11417 13495 11429
rect 13437 11383 13449 11417
rect 13483 11383 13495 11417
rect 13437 11371 13495 11383
rect 12893 11005 12951 11017
rect 13464 11006 13492 11371
rect 12893 10971 12905 11005
rect 12939 10971 12951 11005
rect 12893 10959 12951 10971
rect 13448 10994 13508 11006
rect 12908 10780 12936 10959
rect 13448 10942 13450 10994
rect 13502 10942 13508 10994
rect 13448 10925 13508 10942
rect 13448 10891 13461 10925
rect 13495 10891 13508 10925
rect 13448 10878 13508 10891
rect 12774 10766 13044 10780
rect 12774 10526 12780 10766
rect 13020 10526 13044 10766
rect 12774 10510 13044 10526
rect 13616 10449 13644 12118
rect 13940 12078 13968 12118
rect 13924 12065 13986 12078
rect 13924 12031 13937 12065
rect 13971 12031 13986 12065
rect 13924 12018 13986 12031
rect 14733 12069 14791 12081
rect 14733 12035 14745 12069
rect 14779 12066 14791 12069
rect 15190 12066 15218 13158
rect 15287 13155 15299 13158
rect 15333 13155 15345 13189
rect 15827 13193 15839 13227
rect 15873 13193 15885 13227
rect 15827 13181 15885 13193
rect 15287 13143 15345 13155
rect 15282 13032 15350 13038
rect 15282 12980 15290 13032
rect 15342 12980 15350 13032
rect 15282 12974 15350 12980
rect 15286 12866 15436 12878
rect 15286 12857 15372 12866
rect 15286 12823 15299 12857
rect 15333 12823 15372 12857
rect 15286 12814 15372 12823
rect 15424 12814 15436 12866
rect 15286 12802 15436 12814
rect 15842 12812 15870 13181
rect 16394 13159 16422 13490
rect 16920 13374 16948 13572
rect 16814 13346 16948 13374
rect 16391 13147 16449 13159
rect 16391 13113 16403 13147
rect 16437 13113 16449 13147
rect 16391 13101 16449 13113
rect 16259 12824 16333 12835
rect 16259 12812 16270 12824
rect 15842 12784 16270 12812
rect 15842 12747 15870 12784
rect 16259 12772 16270 12784
rect 16322 12772 16333 12824
rect 16259 12761 16333 12772
rect 15827 12735 15885 12747
rect 15827 12701 15839 12735
rect 15873 12701 15885 12735
rect 15827 12689 15885 12701
rect 15927 12744 16001 12755
rect 15927 12692 15938 12744
rect 15990 12692 16001 12744
rect 15927 12681 16001 12692
rect 14779 12038 15218 12066
rect 14779 12035 14791 12038
rect 14733 12023 14791 12035
rect 13940 11986 13968 12018
rect 14033 11989 14091 12001
rect 14033 11986 14045 11989
rect 13940 11958 14045 11986
rect 13940 11585 13968 11958
rect 14033 11955 14045 11958
rect 14079 11986 14091 11989
rect 14136 11989 14198 12002
rect 14136 11986 14149 11989
rect 14079 11958 14149 11986
rect 14079 11955 14091 11958
rect 14033 11943 14091 11955
rect 14136 11955 14149 11958
rect 14183 11986 14198 11989
rect 14629 11998 14703 12009
rect 14629 11986 14640 11998
rect 14183 11958 14640 11986
rect 14183 11955 14198 11958
rect 14136 11942 14198 11955
rect 14260 11921 14288 11958
rect 14629 11946 14640 11958
rect 14692 11946 14703 11998
rect 14629 11935 14703 11946
rect 14245 11909 14303 11921
rect 14245 11875 14257 11909
rect 14291 11875 14303 11909
rect 14245 11863 14303 11875
rect 14748 11589 14776 12023
rect 15297 11989 15355 12001
rect 15297 11955 15309 11989
rect 15343 11955 15355 11989
rect 15297 11943 15355 11955
rect 15861 11989 15919 12001
rect 15861 11955 15873 11989
rect 15907 11955 15919 11989
rect 15861 11943 15919 11955
rect 13925 11573 13983 11585
rect 13925 11539 13937 11573
rect 13971 11539 13983 11573
rect 13925 11527 13983 11539
rect 14733 11577 14791 11589
rect 14733 11543 14745 11577
rect 14779 11543 14791 11577
rect 14733 11531 14791 11543
rect 13940 11494 13968 11527
rect 14033 11497 14091 11509
rect 14033 11494 14045 11497
rect 13940 11466 14045 11494
rect 14033 11463 14045 11466
rect 14079 11494 14091 11497
rect 14137 11497 14195 11509
rect 14137 11494 14149 11497
rect 14079 11466 14149 11494
rect 14079 11463 14091 11466
rect 14033 11451 14091 11463
rect 14137 11463 14149 11466
rect 14183 11463 14195 11497
rect 14137 11451 14195 11463
rect 13927 11426 14001 11437
rect 13927 11374 13938 11426
rect 13990 11374 14001 11426
rect 14152 11414 14180 11451
rect 14245 11417 14303 11429
rect 14245 11414 14257 11417
rect 14152 11386 14257 11414
rect 13927 11363 14001 11374
rect 14245 11383 14257 11386
rect 14291 11383 14303 11417
rect 14245 11371 14303 11383
rect 13950 11108 13978 11363
rect 13858 11081 14314 11108
rect 14748 11097 14776 11531
rect 15312 11509 15340 11943
rect 15878 11509 15906 11943
rect 15950 11906 15978 12681
rect 16406 12667 16434 13101
rect 16391 12655 16449 12667
rect 16391 12621 16403 12655
rect 16437 12621 16449 12655
rect 16391 12609 16449 12621
rect 16814 12064 16842 13346
rect 17702 13319 17730 13753
rect 18146 13734 18154 13947
rect 18367 13734 18382 13947
rect 18146 13719 18382 13734
rect 18146 13685 18243 13719
rect 18277 13685 18382 13719
rect 18146 13668 18382 13685
rect 16879 13305 16937 13317
rect 16879 13271 16891 13305
rect 16925 13302 16937 13305
rect 17687 13307 17745 13319
rect 16925 13274 17030 13302
rect 16925 13271 16937 13274
rect 16879 13259 16937 13271
rect 17002 13239 17030 13274
rect 17687 13273 17699 13307
rect 17733 13273 17745 13307
rect 17687 13261 17745 13273
rect 16987 13227 17045 13239
rect 16987 13193 16999 13227
rect 17033 13224 17045 13227
rect 17091 13227 17149 13239
rect 17091 13224 17103 13227
rect 17033 13196 17103 13224
rect 17033 13193 17045 13196
rect 16987 13181 17045 13193
rect 17091 13193 17103 13196
rect 17137 13224 17149 13227
rect 17137 13196 17242 13224
rect 17137 13193 17149 13196
rect 17091 13181 17149 13193
rect 17214 13161 17242 13196
rect 17199 13149 17257 13161
rect 17199 13146 17211 13149
rect 17122 13118 17211 13146
rect 16879 12813 16937 12825
rect 16879 12779 16891 12813
rect 16925 12779 16937 12813
rect 16879 12767 16937 12779
rect 16894 12732 16922 12767
rect 17122 12747 17150 13118
rect 17199 13115 17211 13118
rect 17245 13115 17257 13149
rect 17199 13103 17257 13115
rect 17179 12824 17253 12835
rect 17702 12827 17730 13261
rect 18246 13239 18274 13668
rect 18391 13556 18465 13567
rect 18391 13504 18402 13556
rect 18454 13544 18465 13556
rect 19022 13544 19050 13995
rect 19218 13647 19246 14010
rect 19769 13996 19780 14010
rect 19832 13996 19843 14048
rect 19769 13985 19843 13996
rect 20546 13854 20598 13860
rect 20546 13796 20598 13802
rect 19195 13636 19269 13647
rect 19195 13584 19206 13636
rect 19258 13584 19269 13636
rect 19195 13573 19269 13584
rect 18454 13516 19908 13544
rect 18454 13504 18465 13516
rect 18391 13493 18465 13504
rect 19087 13474 19161 13485
rect 19087 13422 19098 13474
rect 19150 13450 19161 13474
rect 19194 13474 19270 13486
rect 19194 13450 19206 13474
rect 19150 13422 19206 13450
rect 19258 13422 19270 13474
rect 19880 13463 19908 13516
rect 19087 13419 19107 13422
rect 19141 13419 19161 13422
rect 19087 13411 19161 13419
rect 19095 13407 19153 13411
rect 19194 13410 19270 13422
rect 19865 13451 19923 13463
rect 19865 13417 19877 13451
rect 19911 13448 19923 13451
rect 19911 13420 20016 13448
rect 19911 13417 19923 13420
rect 18853 13373 18911 13385
rect 18853 13339 18865 13373
rect 18899 13370 18911 13373
rect 19101 13370 19175 13375
rect 18899 13364 19175 13370
rect 18899 13342 19112 13364
rect 18899 13339 18911 13342
rect 18853 13327 18911 13339
rect 18246 13227 18309 13239
rect 18246 13196 18263 13227
rect 18251 13193 18263 13196
rect 18297 13193 18309 13227
rect 18251 13181 18309 13193
rect 18952 13218 18980 13342
rect 19101 13312 19112 13342
rect 19164 13312 19175 13364
rect 19208 13373 19262 13410
rect 19865 13405 19923 13417
rect 19988 13385 20016 13420
rect 19413 13375 19471 13385
rect 19208 13339 19215 13373
rect 19249 13339 19262 13373
rect 19208 13326 19262 13339
rect 19405 13373 19479 13375
rect 19405 13364 19425 13373
rect 19459 13364 19479 13373
rect 19009 13293 19067 13305
rect 19101 13301 19175 13312
rect 19405 13312 19416 13364
rect 19468 13312 19479 13364
rect 19973 13373 20031 13385
rect 19973 13339 19985 13373
rect 20019 13339 20031 13373
rect 19973 13327 20031 13339
rect 19405 13301 19479 13312
rect 19009 13259 19021 13293
rect 19055 13272 19067 13293
rect 19677 13293 19735 13305
rect 19677 13272 19689 13293
rect 19055 13259 19689 13272
rect 19723 13259 19735 13293
rect 19009 13247 19735 13259
rect 19024 13244 19720 13247
rect 18952 13190 18988 13218
rect 18163 13140 18237 13151
rect 18163 13088 18174 13140
rect 18226 13088 18237 13140
rect 18163 13077 18237 13088
rect 17179 12772 17190 12824
rect 17242 12812 17253 12824
rect 17687 12815 17745 12827
rect 17687 12812 17699 12815
rect 17242 12784 17699 12812
rect 17242 12772 17253 12784
rect 17179 12761 17253 12772
rect 17687 12781 17699 12784
rect 17733 12781 17745 12815
rect 17687 12769 17745 12781
rect 16987 12735 17045 12747
rect 16987 12732 16999 12735
rect 16894 12704 16999 12732
rect 16987 12701 16999 12704
rect 17033 12732 17045 12735
rect 17091 12735 17150 12747
rect 17091 12732 17103 12735
rect 17033 12704 17103 12732
rect 17033 12701 17045 12704
rect 16987 12689 17045 12701
rect 17091 12701 17103 12704
rect 17137 12732 17150 12735
rect 18186 12732 18214 13077
rect 18266 12747 18294 13181
rect 18857 13084 18931 13095
rect 18857 13072 18868 13084
rect 18798 13044 18868 13072
rect 18798 12886 18826 13044
rect 18857 13032 18868 13044
rect 18920 13032 18931 13084
rect 18857 13021 18931 13032
rect 18857 12978 18931 12989
rect 18857 12926 18868 12978
rect 18920 12926 18931 12978
rect 18857 12915 18931 12926
rect 18798 12858 18874 12886
rect 17137 12704 18214 12732
rect 18251 12735 18309 12747
rect 17137 12701 17149 12704
rect 17091 12689 17149 12701
rect 16898 12067 16974 12088
rect 16898 12064 16917 12067
rect 16814 12036 16917 12064
rect 16898 12033 16917 12036
rect 16951 12033 16974 12067
rect 17002 12066 17030 12689
rect 17214 12669 17242 12704
rect 18251 12701 18263 12735
rect 18297 12701 18309 12735
rect 18251 12689 18309 12701
rect 17199 12657 17257 12669
rect 17199 12623 17211 12657
rect 17245 12623 17257 12657
rect 17199 12611 17257 12623
rect 17205 12078 17279 12089
rect 17205 12066 17216 12078
rect 17002 12038 17216 12066
rect 16898 12012 16974 12033
rect 17205 12026 17216 12038
rect 17268 12026 17279 12078
rect 17205 12015 17279 12026
rect 17711 12069 17769 12081
rect 17711 12035 17723 12069
rect 17757 12035 17769 12069
rect 17711 12023 17769 12035
rect 16920 12002 16974 12012
rect 16920 11989 17176 12002
rect 16920 11955 17023 11989
rect 17057 11955 17129 11989
rect 17163 11986 17176 11989
rect 17163 11974 17362 11986
rect 17163 11955 17298 11974
rect 16920 11936 17298 11955
rect 16993 11935 17067 11936
rect 17224 11922 17298 11936
rect 17350 11922 17362 11974
rect 16417 11909 16475 11921
rect 16417 11906 16429 11909
rect 15950 11878 16429 11906
rect 16417 11875 16429 11878
rect 16463 11875 16475 11909
rect 16417 11863 16475 11875
rect 17224 11911 17362 11922
rect 17224 11877 17237 11911
rect 17271 11877 17362 11911
rect 17224 11864 17362 11877
rect 15297 11497 15355 11509
rect 15297 11463 15309 11497
rect 15343 11463 15355 11497
rect 15297 11451 15355 11463
rect 15863 11497 15921 11509
rect 15863 11463 15875 11497
rect 15909 11463 15921 11497
rect 15863 11451 15921 11463
rect 13858 11047 13947 11081
rect 13981 11047 14314 11081
rect 13858 11005 14314 11047
rect 14743 11085 14801 11097
rect 14743 11051 14755 11085
rect 14789 11051 14801 11085
rect 14743 11039 14801 11051
rect 15312 11017 15340 11451
rect 15878 11082 15906 11451
rect 16432 11429 16460 11863
rect 17205 11666 17279 11677
rect 17205 11654 17216 11666
rect 17002 11626 17216 11654
rect 16915 11575 16973 11587
rect 16915 11541 16927 11575
rect 16961 11572 16973 11575
rect 17002 11572 17030 11626
rect 17205 11614 17216 11626
rect 17268 11614 17279 11666
rect 17205 11603 17279 11614
rect 17738 11589 17766 12023
rect 18267 11989 18325 12001
rect 18267 11986 18279 11989
rect 17818 11985 18279 11986
rect 17795 11974 18279 11985
rect 17795 11922 17806 11974
rect 17858 11958 18279 11974
rect 17858 11922 17869 11958
rect 18267 11955 18279 11958
rect 18313 11986 18325 11989
rect 18846 11986 18874 12858
rect 18313 11958 18874 11986
rect 18960 12867 18988 13190
rect 19051 13198 19125 13209
rect 19051 13146 19062 13198
rect 19114 13146 19125 13198
rect 19051 13135 19125 13146
rect 19349 13164 19423 13175
rect 19074 13094 19102 13135
rect 19349 13112 19360 13164
rect 19412 13112 19423 13164
rect 19349 13101 19423 13112
rect 19056 13084 19120 13094
rect 19056 13032 19062 13084
rect 19114 13032 19120 13084
rect 19056 13022 19120 13032
rect 19071 12978 19145 12989
rect 19372 12987 19400 13101
rect 19071 12926 19082 12978
rect 19134 12966 19145 12978
rect 19349 12976 19423 12987
rect 19349 12966 19360 12976
rect 19134 12938 19360 12966
rect 19134 12926 19145 12938
rect 19071 12915 19145 12926
rect 19349 12924 19360 12938
rect 19412 12924 19423 12976
rect 19349 12913 19423 12924
rect 18960 12861 19091 12867
rect 18960 12740 18970 12861
rect 19091 12786 19092 12814
rect 18960 12734 19091 12740
rect 18313 11955 18330 11958
rect 18267 11943 18330 11955
rect 17795 11911 17869 11922
rect 17723 11577 17781 11589
rect 16961 11544 17066 11572
rect 16961 11541 16973 11544
rect 16915 11529 16973 11541
rect 17038 11509 17066 11544
rect 17723 11543 17735 11577
rect 17769 11543 17781 11577
rect 17723 11531 17781 11543
rect 17023 11497 17081 11509
rect 17023 11463 17035 11497
rect 17069 11494 17081 11497
rect 17127 11497 17185 11509
rect 17127 11494 17139 11497
rect 17069 11466 17139 11494
rect 17069 11463 17081 11466
rect 17023 11451 17081 11463
rect 17127 11463 17139 11466
rect 17173 11494 17185 11497
rect 17173 11466 17278 11494
rect 17173 11463 17185 11466
rect 17127 11451 17185 11463
rect 17250 11431 17278 11466
rect 16427 11417 16485 11429
rect 16427 11383 16439 11417
rect 16473 11383 16485 11417
rect 17235 11419 17293 11431
rect 17235 11416 17247 11419
rect 16427 11371 16485 11383
rect 17160 11388 17247 11416
rect 16442 11185 16470 11371
rect 16419 11174 16493 11185
rect 16419 11122 16430 11174
rect 16482 11122 16493 11174
rect 16419 11111 16493 11122
rect 16789 11094 16863 11105
rect 16789 11082 16800 11094
rect 15878 11054 16800 11082
rect 15878 11017 15906 11054
rect 16789 11042 16800 11054
rect 16852 11042 16863 11094
rect 16789 11031 16863 11042
rect 16915 11083 16973 11095
rect 16915 11049 16927 11083
rect 16961 11049 16973 11083
rect 16915 11037 16973 11049
rect 15299 11005 15357 11017
rect 13858 10971 14055 11005
rect 14089 10971 14161 11005
rect 14195 10971 14314 11005
rect 13858 10925 14314 10971
rect 14567 10994 14641 11005
rect 14567 10942 14578 10994
rect 14630 10982 14641 10994
rect 15299 10982 15311 11005
rect 14630 10971 15311 10982
rect 15345 10971 15357 11005
rect 14630 10959 15357 10971
rect 15863 11005 15921 11017
rect 15863 10971 15875 11005
rect 15909 10971 15921 11005
rect 15863 10959 15921 10971
rect 16418 11014 16494 11026
rect 16418 10962 16430 11014
rect 16482 10962 16494 11014
rect 16930 11002 16958 11037
rect 17160 11018 17188 11388
rect 17235 11385 17247 11388
rect 17281 11385 17293 11419
rect 17235 11373 17293 11385
rect 17217 11094 17291 11105
rect 17738 11097 17766 11531
rect 18302 11509 18330 11943
rect 18287 11497 18345 11509
rect 18287 11463 18299 11497
rect 18333 11463 18345 11497
rect 18287 11451 18345 11463
rect 17217 11042 17228 11094
rect 17280 11082 17291 11094
rect 17723 11085 17781 11097
rect 17723 11082 17735 11085
rect 17280 11054 17735 11082
rect 17280 11042 17291 11054
rect 17217 11031 17291 11042
rect 17723 11051 17735 11054
rect 17769 11051 17781 11085
rect 17723 11039 17781 11051
rect 17022 11005 17188 11018
rect 18302 11017 18330 11451
rect 17022 11002 17035 11005
rect 16930 10974 17035 11002
rect 14630 10954 15340 10959
rect 14630 10942 14641 10954
rect 14567 10931 14641 10942
rect 13858 10891 14267 10925
rect 14301 10891 14314 10925
rect 13858 10878 14314 10891
rect 16418 10925 16494 10962
rect 17022 10971 17035 10974
rect 17069 10971 17139 11005
rect 17173 10971 17188 11005
rect 17022 10956 17188 10971
rect 18287 11005 18345 11017
rect 18287 10971 18299 11005
rect 18333 10971 18345 11005
rect 18287 10959 18345 10971
rect 16418 10891 16439 10925
rect 16473 10891 16494 10925
rect 16418 10882 16494 10891
rect 17128 10927 17296 10956
rect 18960 10937 18988 12734
rect 19025 11981 19083 11993
rect 19025 11947 19037 11981
rect 19071 11978 19083 11981
rect 19349 11990 19423 12001
rect 19349 11978 19360 11990
rect 19071 11950 19360 11978
rect 19071 11947 19083 11950
rect 19025 11935 19083 11947
rect 19349 11938 19360 11950
rect 19412 11938 19423 11990
rect 17128 10893 17247 10927
rect 17281 10893 17296 10927
rect 17128 10878 17296 10893
rect 18945 10925 19003 10937
rect 18945 10891 18957 10925
rect 18991 10891 19003 10925
rect 18945 10879 19003 10891
rect 13593 10438 13667 10449
rect 13593 10386 13604 10438
rect 13656 10386 13667 10438
rect 13593 10375 13667 10386
rect 13217 10349 13275 10361
rect 13217 10315 13229 10349
rect 13263 10346 13275 10349
rect 13709 10349 13767 10361
rect 13709 10346 13721 10349
rect 13263 10318 13721 10346
rect 13263 10315 13275 10318
rect 13217 10303 13275 10315
rect 13137 9285 13195 9297
rect 13137 9251 13149 9285
rect 13183 9282 13195 9285
rect 13369 9294 13443 9305
rect 13369 9282 13380 9294
rect 13183 9254 13380 9282
rect 13183 9251 13195 9254
rect 13137 9239 13195 9251
rect 13369 9242 13380 9254
rect 13432 9242 13443 9294
rect 13369 9231 13443 9242
rect 13288 8306 13356 8314
rect 13288 8254 13294 8306
rect 13346 8254 13356 8306
rect 13288 8246 13356 8254
rect 13103 8189 13161 8201
rect 13103 8155 13115 8189
rect 13149 8186 13161 8189
rect 13369 8198 13443 8209
rect 13369 8186 13380 8198
rect 13149 8158 13380 8186
rect 13149 8155 13161 8158
rect 13103 8143 13161 8155
rect 13369 8146 13380 8158
rect 13432 8146 13443 8198
rect 13118 7902 13146 8143
rect 13369 8135 13443 8146
rect 13484 7981 13512 10318
rect 13709 10315 13721 10318
rect 13755 10315 13767 10349
rect 13709 10303 13767 10315
rect 13860 9381 13888 10878
rect 19040 10850 19068 11935
rect 19349 11927 19423 11938
rect 19452 10927 19480 13244
rect 19988 13090 20016 13327
rect 19551 13075 19609 13087
rect 19551 13041 19563 13075
rect 19597 13072 19609 13075
rect 19988 13075 20102 13090
rect 19988 13072 20055 13075
rect 19597 13044 20055 13072
rect 19597 13041 19609 13044
rect 19551 13029 19609 13041
rect 20016 13041 20055 13044
rect 20089 13041 20102 13075
rect 20016 13026 20102 13041
rect 19843 12976 19917 12987
rect 19843 12924 19854 12976
rect 19906 12924 19917 12976
rect 19843 12913 19917 12924
rect 19910 12082 20178 12100
rect 19509 11990 19583 12001
rect 19509 11938 19520 11990
rect 19572 11976 19583 11990
rect 19910 11976 19922 12082
rect 19572 11948 19922 11976
rect 19572 11938 19583 11948
rect 19509 11927 19583 11938
rect 19910 11842 19922 11948
rect 20162 11842 20178 12082
rect 19910 11820 20178 11842
rect 19437 10915 19495 10927
rect 19437 10881 19449 10915
rect 19483 10912 19495 10915
rect 19929 10915 19987 10927
rect 19929 10912 19941 10915
rect 19483 10884 19941 10912
rect 19483 10881 19495 10884
rect 19437 10869 19495 10881
rect 19929 10881 19941 10884
rect 19975 10881 19987 10915
rect 19929 10869 19987 10881
rect 14136 10822 19068 10850
rect 13837 9370 13911 9381
rect 13837 9318 13848 9370
rect 13900 9318 13911 9370
rect 13837 9307 13911 9318
rect 13541 9304 13615 9305
rect 13540 9294 13700 9304
rect 13540 9242 13552 9294
rect 13604 9285 13700 9294
rect 14136 9293 14164 10822
rect 14201 10337 14259 10349
rect 14201 10303 14213 10337
rect 14247 10303 14259 10337
rect 14201 10291 14259 10303
rect 14216 10242 14244 10291
rect 14460 10242 14730 10260
rect 14216 10002 14476 10242
rect 14716 10002 14730 10242
rect 13604 9251 13641 9285
rect 13675 9278 13700 9285
rect 14121 9281 14179 9293
rect 14121 9278 14133 9281
rect 13675 9251 14133 9278
rect 13604 9250 14133 9251
rect 13604 9242 13700 9250
rect 13540 9230 13700 9242
rect 14121 9247 14133 9250
rect 14167 9247 14179 9281
rect 14121 9235 14179 9247
rect 13541 8306 13615 8317
rect 13541 8254 13552 8306
rect 13604 8294 13615 8306
rect 13787 8297 13845 8309
rect 13787 8294 13799 8297
rect 13604 8266 13799 8294
rect 13604 8254 13615 8266
rect 13541 8243 13615 8254
rect 13787 8263 13799 8266
rect 13833 8292 13845 8297
rect 14049 8304 14123 8315
rect 14049 8292 14060 8304
rect 13833 8264 14060 8292
rect 13833 8263 13845 8264
rect 13787 8251 13845 8263
rect 14049 8252 14060 8264
rect 14112 8252 14123 8304
rect 14049 8241 14123 8252
rect 13590 8198 13660 8204
rect 13590 8146 13600 8198
rect 13652 8146 13660 8198
rect 13590 8136 13660 8146
rect 13837 8198 13911 8209
rect 13837 8146 13848 8198
rect 13900 8186 13911 8198
rect 14087 8189 14145 8201
rect 14087 8186 14099 8189
rect 13900 8158 14099 8186
rect 13900 8146 13911 8158
rect 13837 8135 13911 8146
rect 14087 8155 14099 8158
rect 14133 8155 14145 8189
rect 14087 8144 14145 8155
rect 14216 8038 14244 10002
rect 14460 9980 14730 10002
rect 19062 9470 19340 9482
rect 19058 8916 19068 9470
rect 19334 8916 19344 9470
rect 19062 8904 19340 8916
rect 18145 8827 18203 8839
rect 18145 8793 18157 8827
rect 18191 8793 18203 8827
rect 18145 8781 18203 8793
rect 17051 8747 17109 8759
rect 17051 8713 17063 8747
rect 17097 8744 17109 8747
rect 17097 8716 17202 8744
rect 17097 8713 17109 8716
rect 17051 8701 17109 8713
rect 17174 8679 17202 8716
rect 17159 8667 17217 8679
rect 17159 8664 17171 8667
rect 16982 8636 17171 8664
rect 14273 8304 14347 8315
rect 14273 8252 14284 8304
rect 14336 8298 14347 8304
rect 14336 8270 15004 8298
rect 14336 8252 14347 8270
rect 14273 8241 14347 8252
rect 14216 8010 14256 8038
rect 13469 7969 13527 7981
rect 13469 7935 13481 7969
rect 13515 7966 13527 7969
rect 13631 7978 13705 7989
rect 13631 7966 13642 7978
rect 13515 7938 13642 7966
rect 13515 7935 13527 7938
rect 13469 7923 13527 7935
rect 13631 7926 13642 7938
rect 13694 7926 13705 7978
rect 14087 7981 14161 7989
rect 14087 7978 14195 7981
rect 13631 7915 13705 7926
rect 13748 7930 14058 7958
rect 13118 7889 13232 7902
rect 13748 7901 13776 7930
rect 13118 7858 13185 7889
rect 13173 7855 13185 7858
rect 13219 7858 13232 7889
rect 13733 7889 13791 7901
rect 13219 7855 13231 7858
rect 13173 7843 13231 7855
rect 13733 7855 13745 7889
rect 13779 7855 13791 7889
rect 13733 7843 13791 7855
rect 13942 7889 14002 7902
rect 13942 7855 13955 7889
rect 13989 7855 14002 7889
rect 14030 7886 14058 7930
rect 14087 7926 14098 7978
rect 14150 7969 14195 7978
rect 14183 7935 14195 7969
rect 14150 7926 14195 7935
rect 14087 7923 14195 7926
rect 14087 7915 14161 7923
rect 14228 7886 14256 8010
rect 14293 7889 14351 7901
rect 14293 7886 14305 7889
rect 14030 7858 14305 7886
rect 13188 7810 13216 7843
rect 13942 7830 14002 7855
rect 14293 7855 14305 7858
rect 14339 7855 14351 7889
rect 14293 7843 14351 7855
rect 13281 7813 13339 7825
rect 13281 7810 13293 7813
rect 13188 7782 13293 7810
rect 13281 7779 13293 7782
rect 13327 7779 13339 7813
rect 13281 7767 13339 7779
rect 13942 7811 14108 7830
rect 13942 7777 14061 7811
rect 14095 7777 14108 7811
rect 13296 7174 13324 7767
rect 13942 7764 14108 7777
rect 13978 7662 14030 7764
rect 13978 7604 14030 7610
rect 13867 7255 13925 7267
rect 13867 7221 13879 7255
rect 13913 7252 13925 7255
rect 13990 7252 14018 7604
rect 14976 7347 15004 8270
rect 16982 7680 17010 8636
rect 17159 8633 17171 8636
rect 17205 8633 17217 8667
rect 17159 8621 17217 8633
rect 18160 8347 18188 8781
rect 19201 8747 19259 8759
rect 19201 8713 19213 8747
rect 19247 8713 19259 8747
rect 19201 8701 19259 8713
rect 18135 8335 18193 8347
rect 18135 8301 18147 8335
rect 18181 8301 18193 8335
rect 18135 8289 18193 8301
rect 17039 8255 17097 8267
rect 17039 8221 17051 8255
rect 17085 8252 17097 8255
rect 17085 8224 17190 8252
rect 17085 8221 17097 8224
rect 17039 8209 17097 8221
rect 17162 8187 17190 8224
rect 17147 8175 17205 8187
rect 17147 8141 17159 8175
rect 17193 8141 17205 8175
rect 17147 8129 17205 8141
rect 17039 7763 17097 7775
rect 17039 7729 17051 7763
rect 17085 7760 17097 7763
rect 17162 7760 17190 8129
rect 18150 7855 18178 8289
rect 19216 8267 19244 8701
rect 19199 8255 19257 8267
rect 19199 8221 19211 8255
rect 19245 8221 19257 8255
rect 19199 8209 19257 8221
rect 18135 7843 18193 7855
rect 18135 7809 18147 7843
rect 18181 7809 18193 7843
rect 18135 7797 18193 7809
rect 19214 7775 19242 8209
rect 19199 7763 19257 7775
rect 19199 7760 19211 7763
rect 17085 7732 17190 7760
rect 17085 7729 17097 7732
rect 17039 7717 17097 7729
rect 17162 7695 17190 7732
rect 18224 7732 19211 7760
rect 17147 7683 17205 7695
rect 16982 7652 17078 7680
rect 14961 7335 15019 7347
rect 14961 7301 14973 7335
rect 15007 7301 15019 7335
rect 14961 7289 15019 7301
rect 13913 7224 14018 7252
rect 13913 7221 13925 7224
rect 13867 7209 13925 7221
rect 13990 7189 14018 7224
rect 13975 7177 14033 7189
rect 13296 7146 13898 7174
rect 13870 6775 13898 7146
rect 13975 7143 13987 7177
rect 14021 7148 14033 7177
rect 14841 7160 14915 7171
rect 14841 7148 14852 7160
rect 14021 7143 14852 7148
rect 13975 7131 14852 7143
rect 13990 7120 14852 7131
rect 14841 7108 14852 7120
rect 14904 7108 14915 7160
rect 14841 7097 14915 7108
rect 14976 6855 15004 7289
rect 16017 7255 16075 7267
rect 16017 7221 16029 7255
rect 16063 7221 16075 7255
rect 16017 7209 16075 7221
rect 15033 7160 15107 7171
rect 15033 7108 15044 7160
rect 15096 7148 15107 7160
rect 15927 7160 16001 7171
rect 15927 7148 15938 7160
rect 15096 7120 15938 7148
rect 15096 7108 15107 7120
rect 15033 7097 15107 7108
rect 15927 7108 15938 7120
rect 15990 7108 16001 7160
rect 15927 7097 16001 7108
rect 14951 6843 15009 6855
rect 14951 6809 14963 6843
rect 14997 6809 15009 6843
rect 14951 6797 15009 6809
rect 13855 6763 13913 6775
rect 13855 6729 13867 6763
rect 13901 6760 13913 6763
rect 13901 6732 14006 6760
rect 13901 6729 13913 6732
rect 13855 6717 13913 6729
rect 13870 6283 13898 6717
rect 13978 6697 14006 6732
rect 13963 6685 14021 6697
rect 13963 6651 13975 6685
rect 14009 6651 14021 6685
rect 13963 6639 14021 6651
rect 13855 6271 13913 6283
rect 13855 6237 13867 6271
rect 13901 6268 13913 6271
rect 13978 6268 14006 6639
rect 14966 6363 14994 6797
rect 16032 6775 16060 7209
rect 17050 7174 17078 7652
rect 17147 7649 17159 7683
rect 17193 7649 17205 7683
rect 17147 7637 17205 7649
rect 16112 7171 17078 7174
rect 16089 7160 17078 7171
rect 16089 7108 16100 7160
rect 16152 7146 17078 7160
rect 16152 7108 16163 7146
rect 16089 7097 16163 7108
rect 17050 6775 17078 7146
rect 17160 6980 17188 7637
rect 17144 6967 17246 6980
rect 17144 6933 17157 6967
rect 17191 6933 17246 6967
rect 17144 6920 17246 6933
rect 16015 6763 16073 6775
rect 16015 6729 16027 6763
rect 16061 6729 16073 6763
rect 16015 6717 16073 6729
rect 17027 6764 17101 6775
rect 16030 6512 16058 6717
rect 17027 6712 17038 6764
rect 17090 6712 17101 6764
rect 17027 6701 17101 6712
rect 16569 6515 16627 6527
rect 16569 6512 16581 6515
rect 16030 6484 16581 6512
rect 14951 6351 15009 6363
rect 14951 6317 14963 6351
rect 14997 6317 15009 6351
rect 14951 6305 15009 6317
rect 16030 6283 16058 6484
rect 16569 6481 16581 6484
rect 16615 6512 16627 6515
rect 16615 6484 17174 6512
rect 16615 6481 16627 6484
rect 16569 6469 16627 6481
rect 17027 6444 17101 6455
rect 17027 6392 17038 6444
rect 17090 6392 17101 6444
rect 17146 6411 17174 6484
rect 17027 6381 17101 6392
rect 17131 6399 17189 6411
rect 13901 6240 14006 6268
rect 13901 6237 13913 6240
rect 13855 6225 13913 6237
rect 13870 5848 13898 6225
rect 13978 6205 14006 6240
rect 16015 6271 16073 6283
rect 16015 6237 16027 6271
rect 16061 6237 16073 6271
rect 16015 6225 16073 6237
rect 13963 6193 14021 6205
rect 13963 6159 13975 6193
rect 14009 6159 14021 6193
rect 13963 6147 14021 6159
rect 13050 5434 13060 5848
rect 14898 5434 14908 5848
rect 15119 5603 15177 5615
rect 15119 5569 15131 5603
rect 15165 5600 15177 5603
rect 15477 5605 15535 5617
rect 15477 5600 15489 5605
rect 15165 5572 15489 5600
rect 15165 5569 15177 5572
rect 15119 5557 15177 5569
rect 15477 5571 15489 5572
rect 15523 5571 15535 5605
rect 15477 5559 15535 5571
rect 16339 5459 16397 5471
rect 13395 4623 13453 4635
rect 13395 4589 13407 4623
rect 13441 4620 13453 4623
rect 13441 4592 13776 4620
rect 13441 4589 13453 4592
rect 13395 4577 13453 4589
rect 13714 4575 13776 4592
rect 13992 4587 14020 5434
rect 16339 5425 16351 5459
rect 16385 5425 16397 5459
rect 16339 5413 16397 5425
rect 16251 5144 16325 5155
rect 16251 5132 16262 5144
rect 15598 5104 16262 5132
rect 14655 4634 14713 4635
rect 14654 4623 14713 4634
rect 14654 4589 14667 4623
rect 14701 4589 14713 4623
rect 15598 4595 15626 5104
rect 16251 5092 16262 5104
rect 16314 5092 16325 5144
rect 16251 5081 16325 5092
rect 16354 5072 16382 5413
rect 17072 5072 17100 6381
rect 17131 6365 17143 6399
rect 17177 6365 17189 6399
rect 17131 6353 17189 6365
rect 17146 5819 17174 6353
rect 17218 6268 17246 6920
rect 18224 6847 18252 7732
rect 19199 7729 19211 7732
rect 19245 7729 19257 7763
rect 19199 7717 19257 7729
rect 19197 7095 19255 7107
rect 19197 7061 19209 7095
rect 19243 7061 19255 7095
rect 19197 7049 19255 7061
rect 19212 6964 19240 7049
rect 19305 6967 19363 6979
rect 19305 6964 19317 6967
rect 19204 6936 19317 6964
rect 18209 6835 18267 6847
rect 18209 6801 18221 6835
rect 18255 6801 18267 6835
rect 18209 6789 18267 6801
rect 18224 6528 18252 6789
rect 18160 6515 18252 6528
rect 18160 6481 18173 6515
rect 18207 6481 18252 6515
rect 18160 6468 18252 6481
rect 18176 6371 18204 6468
rect 19204 6375 19232 6936
rect 19305 6933 19317 6936
rect 19351 6933 19363 6967
rect 19305 6921 19363 6933
rect 18153 6360 18227 6371
rect 18153 6308 18164 6360
rect 18216 6308 18227 6360
rect 19189 6363 19247 6375
rect 19189 6329 19201 6363
rect 19235 6329 19247 6363
rect 19189 6317 19247 6329
rect 18153 6297 18227 6308
rect 17218 6267 18204 6268
rect 17218 6255 18219 6267
rect 17218 6240 18173 6255
rect 17145 5807 17203 5819
rect 17145 5773 17157 5807
rect 17191 5773 17203 5807
rect 17145 5761 17203 5773
rect 17146 5161 17174 5761
rect 17304 5539 17332 6240
rect 18161 6221 18173 6240
rect 18207 6252 18219 6255
rect 19204 6252 19232 6317
rect 18207 6224 19232 6252
rect 18207 6221 18219 6224
rect 18161 6209 18219 6221
rect 18176 5588 18204 6209
rect 19204 6047 19232 6224
rect 19197 6035 19255 6047
rect 19197 6001 19209 6035
rect 19243 6001 19255 6035
rect 19197 5989 19255 6001
rect 19212 5804 19240 5989
rect 19305 5807 19363 5819
rect 19305 5804 19317 5807
rect 19212 5776 19317 5804
rect 19305 5773 19317 5776
rect 19351 5773 19363 5807
rect 19305 5761 19363 5773
rect 18176 5575 18268 5588
rect 18176 5544 18221 5575
rect 18208 5541 18221 5544
rect 18255 5541 18268 5575
rect 17281 5528 17355 5539
rect 18208 5528 18268 5541
rect 17281 5476 17292 5528
rect 17344 5476 17355 5528
rect 17281 5465 17355 5476
rect 18153 5264 18227 5275
rect 18153 5212 18164 5264
rect 18216 5212 18227 5264
rect 18153 5201 18227 5212
rect 18176 5200 18204 5201
rect 17131 5155 17189 5161
rect 17131 5149 17243 5155
rect 17131 5115 17143 5149
rect 17177 5144 17243 5149
rect 17177 5115 17180 5144
rect 17131 5103 17180 5115
rect 17169 5092 17180 5103
rect 17232 5092 17243 5144
rect 17169 5081 17243 5092
rect 19189 5111 19247 5123
rect 19189 5077 19201 5111
rect 19235 5077 19247 5111
rect 16354 5044 17136 5072
rect 19189 5065 19247 5077
rect 17094 5020 17136 5044
rect 17094 5005 17158 5020
rect 17094 4971 17109 5005
rect 17143 4971 17158 5005
rect 17094 4958 17158 4971
rect 17112 4896 17140 4958
rect 18161 4899 18219 4911
rect 18161 4896 18173 4899
rect 17112 4868 18173 4896
rect 17112 4803 17140 4868
rect 18161 4865 18173 4868
rect 18207 4896 18219 4899
rect 18207 4868 18440 4896
rect 18207 4865 18219 4868
rect 18161 4853 18219 4865
rect 17281 4828 17355 4839
rect 17112 4791 17191 4803
rect 17112 4757 17145 4791
rect 17179 4757 17191 4791
rect 17281 4776 17292 4828
rect 17344 4776 17355 4828
rect 17281 4765 17355 4776
rect 17112 4745 17191 4757
rect 13714 4541 13729 4575
rect 13763 4572 13776 4575
rect 13834 4572 13840 4584
rect 13763 4544 13840 4572
rect 13763 4541 13776 4544
rect 13714 4528 13776 4541
rect 13834 4532 13840 4544
rect 13892 4532 13898 4584
rect 13977 4575 14035 4587
rect 13977 4541 13989 4575
rect 14023 4572 14035 4575
rect 14654 4577 14713 4589
rect 14978 4584 15036 4590
rect 14654 4572 14698 4577
rect 14023 4544 14698 4572
rect 14023 4541 14035 4544
rect 13977 4529 14035 4541
rect 14978 4532 14984 4584
rect 14978 4529 15036 4532
rect 15333 4575 15391 4587
rect 15333 4541 15345 4575
rect 15379 4541 15391 4575
rect 15333 4529 15391 4541
rect 15575 4584 15649 4595
rect 15575 4532 15586 4584
rect 15638 4532 15649 4584
rect 13707 3634 13781 3645
rect 13707 3614 13718 3634
rect 13258 3586 13718 3614
rect 13258 3559 13324 3586
rect 13707 3582 13718 3586
rect 13770 3614 13781 3634
rect 13992 3614 14020 4529
rect 14984 4526 15036 4529
rect 14763 4376 14837 4387
rect 14763 4324 14774 4376
rect 14826 4364 14837 4376
rect 15348 4364 15376 4529
rect 15575 4521 15649 4532
rect 16796 4473 16856 4486
rect 16796 4439 16809 4473
rect 16843 4439 16856 4473
rect 16796 4426 16856 4439
rect 16569 4367 16627 4379
rect 16569 4364 16581 4367
rect 14826 4336 16581 4364
rect 14826 4324 14837 4336
rect 14763 4313 14837 4324
rect 13770 3586 14020 3614
rect 13770 3582 13781 3586
rect 13707 3571 13781 3582
rect 13258 3525 13277 3559
rect 13311 3525 13324 3559
rect 14425 3559 14483 3571
rect 13831 3545 13889 3557
rect 13831 3542 13843 3545
rect 13258 3506 13324 3525
rect 13730 3514 13843 3542
rect 13730 2995 13758 3514
rect 13831 3511 13843 3514
rect 13877 3542 13889 3545
rect 14425 3542 14437 3559
rect 13877 3525 14437 3542
rect 14471 3542 14483 3559
rect 15083 3545 15141 3557
rect 15083 3542 15095 3545
rect 14471 3525 15095 3542
rect 13877 3514 15095 3525
rect 13877 3511 13889 3514
rect 14425 3513 14483 3514
rect 13831 3499 13889 3511
rect 15083 3511 15095 3514
rect 15129 3511 15141 3545
rect 15348 3544 15376 4336
rect 16569 4333 16581 4336
rect 16615 4364 16627 4367
rect 16812 4364 16840 4426
rect 17112 4364 17140 4745
rect 16615 4336 17140 4364
rect 16615 4333 16627 4336
rect 16569 4321 16627 4333
rect 16339 3871 16397 3883
rect 16339 3837 16351 3871
rect 16385 3837 16397 3871
rect 16339 3825 16397 3837
rect 15439 3547 15497 3559
rect 15439 3544 15451 3547
rect 15242 3523 15451 3544
rect 15083 3499 15141 3511
rect 15227 3516 15451 3523
rect 15227 3511 15285 3516
rect 14763 3300 14837 3311
rect 14763 3248 14774 3300
rect 14826 3248 14837 3300
rect 14763 3237 14837 3248
rect 13715 2983 13773 2995
rect 13715 2949 13727 2983
rect 13761 2949 13773 2983
rect 13715 2937 13773 2949
rect 13707 2760 13781 2771
rect 14786 2765 14814 3237
rect 15098 3151 15126 3499
rect 15227 3477 15239 3511
rect 15273 3477 15285 3511
rect 15439 3513 15451 3516
rect 15485 3544 15497 3547
rect 15485 3516 15802 3544
rect 16356 3527 16384 3825
rect 15485 3513 15497 3516
rect 15439 3501 15497 3513
rect 15227 3465 15285 3477
rect 15075 3140 15149 3151
rect 15075 3088 15086 3140
rect 15138 3088 15149 3140
rect 15075 3077 15149 3088
rect 13707 2708 13718 2760
rect 13770 2708 13781 2760
rect 14771 2753 14829 2765
rect 14771 2750 14783 2753
rect 13707 2697 13781 2708
rect 13842 2722 14783 2750
rect 13730 2588 13758 2697
rect 13842 2691 13870 2722
rect 14771 2719 14783 2722
rect 14817 2750 14829 2753
rect 15242 2750 15270 3465
rect 15774 3223 15802 3516
rect 16341 3515 16399 3527
rect 16341 3481 16353 3515
rect 16387 3481 16399 3515
rect 16341 3469 16399 3481
rect 15759 3211 15817 3223
rect 15759 3177 15771 3211
rect 15805 3177 15817 3211
rect 17304 3208 17332 4765
rect 18154 4662 18226 4664
rect 18153 4660 18226 4662
rect 18153 4658 18227 4660
rect 18153 4606 18164 4658
rect 18216 4606 18227 4658
rect 18153 4595 18227 4606
rect 18412 4150 18440 4868
rect 19204 4767 19232 5065
rect 19191 4755 19249 4767
rect 19191 4721 19203 4755
rect 19237 4721 19249 4755
rect 19191 4709 19249 4721
rect 18961 4259 19019 4271
rect 18961 4256 18973 4259
rect 18748 4228 18973 4256
rect 18748 4165 18776 4228
rect 18961 4225 18973 4228
rect 19007 4225 19019 4259
rect 18961 4213 19019 4225
rect 18733 4153 18791 4165
rect 18733 4150 18745 4153
rect 18412 4122 18745 4150
rect 17361 3986 17435 3997
rect 17361 3934 17372 3986
rect 17424 3934 17435 3986
rect 17361 3923 17435 3934
rect 18412 3847 18440 4122
rect 18733 4119 18745 4122
rect 18779 4119 18791 4153
rect 18733 4107 18791 4119
rect 18397 3835 18455 3847
rect 18397 3801 18409 3835
rect 18443 3801 18455 3835
rect 18397 3789 18455 3801
rect 17369 3727 17427 3739
rect 17369 3693 17381 3727
rect 17415 3724 17427 3727
rect 18412 3724 18440 3789
rect 17415 3696 18440 3724
rect 17415 3693 17427 3696
rect 17369 3681 17427 3693
rect 18153 3656 18227 3667
rect 17361 3638 17435 3649
rect 17361 3586 17372 3638
rect 17424 3586 17435 3638
rect 18153 3604 18164 3656
rect 18216 3604 18227 3656
rect 18153 3593 18227 3604
rect 18412 3634 18440 3696
rect 18412 3621 18492 3634
rect 17361 3575 17435 3586
rect 17384 3383 17412 3575
rect 18176 3544 18204 3593
rect 18412 3587 18445 3621
rect 18479 3618 18492 3621
rect 19036 3618 19046 3698
rect 18479 3590 19046 3618
rect 18479 3587 18492 3590
rect 18412 3574 18492 3587
rect 18176 3516 18458 3544
rect 18398 3477 18458 3516
rect 18398 3443 18411 3477
rect 18445 3443 18458 3477
rect 18398 3430 18458 3443
rect 17369 3376 17427 3383
rect 17369 3330 17372 3376
rect 17424 3330 17427 3376
rect 17372 3318 17424 3324
rect 17304 3180 17338 3208
rect 15759 3165 15817 3177
rect 15774 2980 15802 3165
rect 17310 3063 17338 3180
rect 17310 3051 17379 3063
rect 17310 3048 17333 3051
rect 16356 3020 17333 3048
rect 15865 2983 15923 2995
rect 15865 2980 15877 2983
rect 15774 2952 15877 2980
rect 15865 2949 15877 2952
rect 15911 2949 15923 2983
rect 15865 2937 15923 2949
rect 14817 2722 15270 2750
rect 14817 2719 14829 2722
rect 14771 2707 14829 2719
rect 13819 2680 13893 2691
rect 13819 2628 13830 2680
rect 13882 2628 13893 2680
rect 13819 2617 13893 2628
rect 15075 2682 15149 2693
rect 15075 2630 15086 2682
rect 15138 2630 15149 2682
rect 15075 2619 15149 2630
rect 14897 2600 14971 2611
rect 14897 2588 14908 2600
rect 13730 2560 14908 2588
rect 13730 2531 13758 2560
rect 14897 2548 14908 2560
rect 14960 2548 14971 2600
rect 14897 2537 14971 2548
rect 13707 2520 13781 2531
rect 13707 2468 13718 2520
rect 13770 2468 13781 2520
rect 13707 2457 13781 2468
rect 14707 2421 14765 2433
rect 14707 2387 14719 2421
rect 14753 2387 14765 2421
rect 14707 2375 14765 2387
rect 13613 2341 13671 2353
rect 13613 2307 13625 2341
rect 13659 2307 13671 2341
rect 13613 2295 13671 2307
rect 13628 2260 13656 2295
rect 13721 2263 13779 2275
rect 13721 2260 13733 2263
rect 13628 2232 13733 2260
rect 13721 2229 13733 2232
rect 13767 2260 13779 2263
rect 13819 2272 13893 2283
rect 13819 2260 13830 2272
rect 13767 2232 13830 2260
rect 13767 2229 13779 2232
rect 13721 2217 13779 2229
rect 13819 2220 13830 2232
rect 13882 2220 13893 2272
rect 13819 2209 13893 2220
rect 13707 1938 13781 1949
rect 14722 1941 14750 2375
rect 15098 2338 15126 2619
rect 15183 2600 15257 2611
rect 15183 2548 15194 2600
rect 15246 2588 15257 2600
rect 15982 2588 15992 2848
rect 15246 2560 15992 2588
rect 15246 2548 15257 2560
rect 15183 2537 15257 2548
rect 15982 2388 15992 2560
rect 16168 2588 16178 2848
rect 16225 2819 16283 2831
rect 16225 2785 16237 2819
rect 16271 2785 16283 2819
rect 16225 2773 16283 2785
rect 16240 2588 16268 2773
rect 16356 2603 16384 3020
rect 17321 3017 17333 3020
rect 17367 3017 17379 3051
rect 17321 3005 17379 3017
rect 16333 2591 16391 2603
rect 16333 2588 16345 2591
rect 16168 2560 16345 2588
rect 16168 2388 16178 2560
rect 16333 2557 16345 2560
rect 16379 2557 16391 2591
rect 16333 2545 16391 2557
rect 16356 2368 16384 2545
rect 17336 2390 17364 3005
rect 18414 2831 18442 3430
rect 19036 2968 19046 3590
rect 19726 2968 19736 3698
rect 18385 2819 18443 2831
rect 18385 2785 18397 2819
rect 18431 2785 18443 2819
rect 18385 2773 18443 2785
rect 17336 2371 17430 2390
rect 17336 2368 17381 2371
rect 15763 2341 15821 2353
rect 15763 2338 15775 2341
rect 15098 2310 15775 2338
rect 15763 2307 15775 2310
rect 15809 2307 15821 2341
rect 15763 2295 15821 2307
rect 16356 2340 17381 2368
rect 15778 2108 15806 2295
rect 16356 2275 16384 2340
rect 17360 2337 17381 2340
rect 17415 2337 17430 2371
rect 17360 2320 17430 2337
rect 17361 2278 17435 2289
rect 16341 2263 16399 2275
rect 16341 2229 16353 2263
rect 16387 2229 16399 2263
rect 16341 2217 16399 2229
rect 17361 2226 17372 2278
rect 17424 2226 17435 2278
rect 18414 2239 18442 2773
rect 16251 2120 16325 2131
rect 16251 2108 16262 2120
rect 15778 2080 16262 2108
rect 13707 1886 13718 1938
rect 13770 1886 13781 1938
rect 13707 1875 13781 1886
rect 14697 1929 14755 1941
rect 14697 1895 14709 1929
rect 14743 1895 14755 1929
rect 14697 1883 14755 1895
rect 13601 1849 13659 1861
rect 13601 1815 13613 1849
rect 13647 1846 13659 1849
rect 13730 1846 13758 1875
rect 13647 1818 13758 1846
rect 13647 1815 13659 1818
rect 13601 1803 13659 1815
rect 13724 1783 13752 1818
rect 13709 1771 13767 1783
rect 13709 1737 13721 1771
rect 13755 1737 13767 1771
rect 13709 1725 13767 1737
rect 13601 1357 13659 1369
rect 13601 1323 13613 1357
rect 13647 1354 13659 1357
rect 13724 1354 13752 1725
rect 14712 1449 14740 1883
rect 15778 1861 15806 2080
rect 16251 2068 16262 2080
rect 16314 2068 16325 2120
rect 16251 2057 16325 2068
rect 15761 1849 15819 1861
rect 15761 1815 15773 1849
rect 15807 1815 15819 1849
rect 15761 1803 15819 1815
rect 14697 1437 14755 1449
rect 14697 1403 14709 1437
rect 14743 1403 14755 1437
rect 14697 1391 14755 1403
rect 15776 1369 15804 1803
rect 16225 1659 16283 1671
rect 16225 1625 16237 1659
rect 16271 1656 16283 1659
rect 16356 1656 16384 2217
rect 17361 2215 17435 2226
rect 18399 2227 18457 2239
rect 16413 2120 16487 2131
rect 17384 2130 17412 2215
rect 18399 2193 18411 2227
rect 18445 2193 18457 2227
rect 18399 2181 18457 2193
rect 16413 2068 16424 2120
rect 16476 2108 16487 2120
rect 17360 2111 17430 2130
rect 17360 2108 17381 2111
rect 16476 2080 17381 2108
rect 16476 2068 16487 2080
rect 16413 2057 16487 2068
rect 17336 2077 17381 2080
rect 17415 2077 17430 2111
rect 18414 2108 18442 2181
rect 18961 2111 19019 2123
rect 18961 2108 18973 2111
rect 18414 2080 18973 2108
rect 17336 2060 17430 2077
rect 18961 2077 18973 2080
rect 19007 2077 19019 2111
rect 18961 2065 19019 2077
rect 17336 1803 17364 2060
rect 17321 1791 17379 1803
rect 17321 1757 17333 1791
rect 17367 1757 17379 1791
rect 17321 1745 17379 1757
rect 18290 1780 18562 1800
rect 16271 1628 16384 1656
rect 16271 1625 16283 1628
rect 16225 1613 16283 1625
rect 16348 1543 16376 1628
rect 16333 1531 16391 1543
rect 16333 1497 16345 1531
rect 16379 1497 16391 1531
rect 18290 1540 18306 1780
rect 18546 1540 18562 1780
rect 18290 1514 18562 1540
rect 16333 1485 16391 1497
rect 13647 1326 13752 1354
rect 13647 1323 13659 1326
rect 13601 1311 13659 1323
rect 13724 1291 13752 1326
rect 15761 1357 15819 1369
rect 15761 1323 15773 1357
rect 15807 1323 15819 1357
rect 15761 1311 15819 1323
rect 13709 1279 13767 1291
rect 13709 1245 13721 1279
rect 13755 1245 13767 1279
rect 13709 1233 13767 1245
<< via1 >>
rect 4545 22145 4615 22215
rect 5090 22191 5150 22251
rect 5630 22190 5690 22250
rect 6210 22190 6270 22250
rect 6750 22190 6810 22250
rect 7330 22190 7390 22250
rect 7870 22190 7930 22250
rect 8430 22190 8490 22250
rect 8990 22190 9050 22250
rect 9550 22190 9610 22250
rect 10130 22190 10190 22250
rect 10670 22190 10730 22250
rect 11190 22190 11250 22250
rect 11750 22190 11810 22250
rect 12310 22190 12370 22250
rect 12870 22190 12930 22250
rect 13410 22190 13470 22250
rect 13970 22190 14030 22250
rect 14550 22190 14610 22250
rect 15070 22190 15130 22250
rect 15630 22190 15690 22250
rect 16170 22190 16230 22250
rect 16710 22190 16770 22250
rect 17270 22190 17330 22250
rect 18958 21035 19043 21120
rect 19196 16534 19248 16586
rect 19860 16569 20050 16650
rect 19860 16533 19939 16569
rect 19939 16533 19973 16569
rect 19973 16533 20050 16569
rect 19860 16450 20050 16533
rect 19360 15513 19412 15522
rect 19360 15479 19367 15513
rect 19367 15479 19401 15513
rect 19401 15479 19412 15513
rect 19360 15470 19412 15479
rect 13886 14308 13938 14360
rect 14046 14308 14098 14360
rect 19516 14525 19568 14534
rect 19516 14491 19525 14525
rect 19525 14491 19559 14525
rect 19559 14491 19568 14525
rect 19516 14482 19568 14491
rect 13966 14086 14018 14138
rect 19834 14417 19886 14426
rect 19834 14383 19859 14417
rect 19859 14383 19886 14417
rect 19834 14374 19886 14383
rect 18974 14294 19026 14346
rect 20010 14525 20062 14534
rect 20010 14491 20017 14525
rect 20017 14491 20051 14525
rect 20051 14491 20062 14525
rect 20010 14482 20062 14491
rect 19196 14201 19248 14208
rect 19196 14167 19207 14201
rect 19207 14167 19241 14201
rect 19241 14167 19248 14201
rect 19196 14156 19248 14167
rect 19834 14199 19886 14208
rect 19834 14165 19875 14199
rect 19875 14165 19886 14199
rect 19834 14156 19886 14165
rect 19780 14041 19832 14048
rect 12914 13663 12931 13674
rect 12931 13663 13389 13674
rect 13389 13663 13423 13674
rect 13423 13663 13478 13674
rect 12914 13444 13478 13663
rect 13966 13676 14018 13728
rect 13870 13560 13922 13612
rect 13458 13260 13510 13312
rect 14030 13560 14082 13612
rect 14446 13560 14498 13612
rect 15372 13478 15424 13530
rect 15290 13355 15342 13364
rect 15290 13321 15299 13355
rect 15299 13321 15333 13355
rect 15333 13321 15342 13355
rect 15290 13312 15342 13321
rect 15910 13478 15962 13530
rect 16492 13560 16544 13612
rect 13938 13058 13990 13110
rect 13938 12716 13990 12768
rect 12840 12230 13080 12470
rect 13458 12106 13510 12158
rect 13450 10942 13502 10994
rect 12780 10526 13020 10766
rect 15290 13023 15342 13032
rect 15290 12989 15299 13023
rect 15299 12989 15333 13023
rect 15333 12989 15342 13023
rect 15290 12980 15342 12989
rect 15372 12814 15424 12866
rect 16270 12772 16322 12824
rect 15938 12692 15990 12744
rect 14640 11946 14692 11998
rect 13938 11374 13990 11426
rect 18154 13734 18367 13947
rect 18402 13504 18454 13556
rect 19780 14007 19789 14041
rect 19789 14007 19823 14041
rect 19823 14007 19832 14041
rect 19780 13996 19832 14007
rect 20546 13802 20598 13854
rect 19206 13584 19258 13636
rect 19098 13453 19150 13474
rect 19098 13422 19107 13453
rect 19107 13422 19141 13453
rect 19141 13422 19150 13453
rect 19206 13422 19258 13474
rect 19112 13312 19164 13364
rect 19416 13339 19425 13364
rect 19425 13339 19459 13364
rect 19459 13339 19468 13364
rect 19416 13312 19468 13339
rect 18174 13088 18226 13140
rect 17190 12772 17242 12824
rect 18868 13032 18920 13084
rect 18868 12969 18920 12978
rect 18868 12935 18879 12969
rect 18879 12935 18913 12969
rect 18913 12935 18920 12969
rect 18868 12926 18920 12935
rect 17216 12026 17268 12078
rect 17298 11922 17350 11974
rect 17216 11614 17268 11666
rect 17806 11922 17858 11974
rect 19062 13146 19114 13198
rect 19360 13112 19412 13164
rect 19062 13075 19114 13084
rect 19062 13041 19071 13075
rect 19071 13041 19105 13075
rect 19105 13041 19114 13075
rect 19062 13032 19114 13041
rect 19082 12926 19134 12978
rect 19360 12967 19412 12976
rect 19360 12933 19371 12967
rect 19371 12933 19405 12967
rect 19405 12933 19412 12967
rect 19360 12924 19412 12933
rect 18970 12740 19091 12861
rect 16430 11122 16482 11174
rect 16800 11042 16852 11094
rect 14578 10942 14630 10994
rect 16430 10962 16482 11014
rect 17228 11042 17280 11094
rect 19360 11938 19412 11990
rect 13604 10386 13656 10438
rect 13380 9242 13432 9294
rect 13294 8297 13346 8306
rect 13294 8263 13307 8297
rect 13307 8263 13341 8297
rect 13341 8263 13346 8297
rect 13294 8254 13346 8263
rect 13380 8146 13432 8198
rect 19854 12967 19906 12976
rect 19854 12933 19863 12967
rect 19863 12933 19897 12967
rect 19897 12933 19906 12967
rect 19854 12924 19906 12933
rect 19520 11979 19572 11990
rect 19520 11945 19529 11979
rect 19529 11945 19563 11979
rect 19563 11945 19572 11979
rect 19922 11979 20162 12082
rect 19520 11938 19572 11945
rect 19922 11945 20021 11979
rect 20021 11945 20055 11979
rect 20055 11945 20162 11979
rect 19922 11842 20162 11945
rect 13848 9318 13900 9370
rect 13552 9242 13604 9294
rect 14476 10002 14716 10242
rect 13552 8254 13604 8306
rect 14060 8252 14112 8304
rect 13600 8189 13652 8198
rect 13600 8155 13607 8189
rect 13607 8155 13641 8189
rect 13641 8155 13652 8189
rect 13600 8146 13652 8155
rect 13848 8146 13900 8198
rect 19068 8916 19334 9470
rect 14284 8295 14336 8304
rect 14284 8261 14291 8295
rect 14291 8261 14325 8295
rect 14325 8261 14336 8295
rect 14284 8252 14336 8261
rect 13642 7926 13694 7978
rect 14098 7969 14150 7978
rect 14098 7935 14149 7969
rect 14149 7935 14150 7969
rect 14098 7926 14150 7935
rect 13978 7610 14030 7662
rect 14852 7108 14904 7160
rect 15044 7108 15096 7160
rect 15938 7108 15990 7160
rect 16100 7108 16152 7160
rect 17038 6712 17090 6764
rect 17038 6392 17090 6444
rect 13060 5719 14898 5848
rect 13060 5685 13277 5719
rect 13277 5685 13311 5719
rect 13311 5685 14437 5719
rect 14437 5685 14471 5719
rect 14471 5685 14898 5719
rect 13060 5611 14898 5685
rect 13060 5577 13149 5611
rect 13149 5577 13183 5611
rect 13183 5603 14209 5611
rect 13183 5577 13881 5603
rect 13060 5569 13881 5577
rect 13881 5569 13915 5603
rect 13915 5577 14209 5603
rect 14209 5577 14243 5611
rect 14243 5577 14898 5611
rect 13915 5569 14898 5577
rect 13060 5434 14898 5569
rect 16262 5092 16314 5144
rect 18164 6308 18216 6360
rect 17292 5476 17344 5528
rect 18164 5255 18216 5264
rect 18164 5221 18173 5255
rect 18173 5221 18207 5255
rect 18207 5221 18216 5255
rect 18164 5212 18216 5221
rect 17180 5092 17232 5144
rect 17292 4776 17344 4828
rect 13840 4532 13892 4584
rect 14984 4575 15036 4584
rect 14984 4541 14989 4575
rect 14989 4541 15023 4575
rect 15023 4541 15036 4575
rect 14984 4532 15036 4541
rect 15586 4575 15638 4584
rect 15586 4541 15595 4575
rect 15595 4541 15629 4575
rect 15629 4541 15638 4575
rect 15586 4532 15638 4541
rect 13718 3582 13770 3634
rect 14774 4324 14826 4376
rect 14774 3248 14826 3300
rect 15086 3088 15138 3140
rect 13718 2708 13770 2760
rect 18164 4649 18216 4658
rect 18164 4615 18173 4649
rect 18173 4615 18207 4649
rect 18207 4615 18216 4649
rect 18164 4606 18216 4615
rect 17372 3977 17424 3986
rect 17372 3943 17381 3977
rect 17381 3943 17415 3977
rect 17415 3943 17424 3977
rect 17372 3934 17424 3943
rect 17372 3586 17424 3638
rect 18164 3604 18216 3656
rect 17372 3371 17424 3376
rect 17372 3337 17381 3371
rect 17381 3337 17415 3371
rect 17415 3337 17424 3371
rect 17372 3324 17424 3337
rect 13830 2628 13882 2680
rect 15086 2630 15138 2682
rect 14908 2548 14960 2600
rect 13718 2468 13770 2520
rect 13830 2220 13882 2272
rect 15194 2548 15246 2600
rect 15992 2388 16168 2848
rect 19046 3167 19726 3698
rect 19046 3133 19203 3167
rect 19203 3133 19237 3167
rect 19237 3133 19726 3167
rect 19046 2968 19726 3133
rect 17372 2226 17424 2278
rect 13718 1886 13770 1938
rect 16262 2068 16314 2120
rect 16424 2068 16476 2120
rect 18306 1659 18546 1780
rect 18306 1625 18397 1659
rect 18397 1625 18431 1659
rect 18431 1625 18546 1659
rect 18306 1540 18546 1625
<< metal2 >>
rect 5060 22251 5180 22280
rect 4520 22215 4640 22240
rect 4520 22145 4545 22215
rect 4615 22145 4640 22215
rect 5060 22191 5090 22251
rect 5150 22191 5180 22251
rect 5060 22160 5180 22191
rect 5600 22250 5720 22280
rect 5600 22190 5630 22250
rect 5690 22190 5720 22250
rect 5600 22160 5720 22190
rect 6180 22250 6300 22280
rect 6180 22190 6210 22250
rect 6270 22190 6300 22250
rect 6180 22160 6300 22190
rect 6720 22250 6840 22280
rect 6720 22190 6750 22250
rect 6810 22190 6840 22250
rect 6720 22160 6840 22190
rect 7300 22250 7420 22280
rect 7300 22190 7330 22250
rect 7390 22190 7420 22250
rect 7300 22160 7420 22190
rect 7840 22250 7960 22280
rect 7840 22190 7870 22250
rect 7930 22190 7960 22250
rect 7840 22160 7960 22190
rect 8400 22250 8520 22280
rect 8400 22190 8430 22250
rect 8490 22190 8520 22250
rect 8400 22160 8520 22190
rect 8960 22250 9080 22280
rect 8960 22190 8990 22250
rect 9050 22190 9080 22250
rect 8960 22160 9080 22190
rect 9520 22250 9640 22280
rect 9520 22190 9550 22250
rect 9610 22190 9640 22250
rect 9520 22160 9640 22190
rect 10100 22250 10220 22280
rect 10100 22190 10130 22250
rect 10190 22190 10220 22250
rect 10100 22160 10220 22190
rect 10640 22250 10760 22280
rect 10640 22190 10670 22250
rect 10730 22190 10760 22250
rect 10640 22160 10760 22190
rect 11160 22250 11280 22280
rect 11160 22190 11190 22250
rect 11250 22190 11280 22250
rect 11160 22160 11280 22190
rect 11720 22250 11840 22280
rect 11720 22190 11750 22250
rect 11810 22190 11840 22250
rect 11720 22160 11840 22190
rect 12280 22250 12400 22280
rect 12280 22190 12310 22250
rect 12370 22190 12400 22250
rect 12280 22160 12400 22190
rect 12840 22250 12960 22280
rect 12840 22190 12870 22250
rect 12930 22190 12960 22250
rect 12840 22160 12960 22190
rect 13380 22250 13500 22280
rect 13380 22190 13410 22250
rect 13470 22190 13500 22250
rect 13380 22160 13500 22190
rect 13940 22250 14060 22280
rect 13940 22190 13970 22250
rect 14030 22190 14060 22250
rect 13940 22160 14060 22190
rect 14520 22250 14640 22280
rect 14520 22190 14550 22250
rect 14610 22190 14640 22250
rect 14520 22160 14640 22190
rect 15040 22250 15160 22280
rect 15040 22190 15070 22250
rect 15130 22190 15160 22250
rect 15040 22160 15160 22190
rect 15600 22250 15720 22280
rect 15600 22190 15630 22250
rect 15690 22190 15720 22250
rect 15600 22160 15720 22190
rect 16140 22250 16260 22280
rect 16140 22190 16170 22250
rect 16230 22190 16260 22250
rect 16140 22160 16260 22190
rect 16680 22250 16800 22280
rect 16680 22190 16710 22250
rect 16770 22190 16800 22250
rect 16680 22160 16800 22190
rect 17240 22250 17360 22280
rect 17240 22190 17270 22250
rect 17330 22190 17360 22250
rect 17240 22160 17360 22190
rect 4520 22120 4640 22145
rect 22978 21780 23221 21781
rect 22420 21775 22660 21780
rect 22978 21775 23222 21780
rect 24070 21776 24310 21780
rect 24070 21775 24316 21776
rect 24630 21775 24870 21780
rect 25166 21779 25414 21784
rect 25702 21782 25956 21787
rect 21920 21768 22145 21773
rect 21916 21553 21925 21768
rect 22140 21553 22149 21768
rect 18958 21120 19043 21126
rect 18958 20732 19043 21035
rect 18958 20722 20700 20732
rect 18958 16846 18992 20722
rect 18958 16836 20700 16846
rect 13875 14360 13949 14371
rect 13875 14308 13886 14360
rect 13938 14348 13949 14360
rect 14035 14360 14109 14371
rect 14035 14348 14046 14360
rect 13938 14320 14046 14348
rect 13938 14308 13949 14320
rect 13875 14297 13949 14308
rect 14035 14308 14046 14320
rect 14098 14308 14109 14360
rect 14035 14297 14109 14308
rect 18958 14346 19043 16836
rect 19838 16650 20070 16672
rect 19196 16586 19248 16592
rect 19196 16528 19248 16534
rect 18958 14294 18974 14346
rect 19026 14294 19043 14346
rect 18958 14278 19043 14294
rect 19208 14222 19236 16528
rect 19838 16450 19860 16650
rect 20050 16450 20070 16650
rect 19838 16430 20070 16450
rect 19346 15524 19427 15537
rect 19346 15468 19358 15524
rect 19414 15468 19427 15524
rect 19346 15455 19427 15468
rect 19505 14534 19579 14545
rect 19505 14482 19516 14534
rect 19568 14522 19579 14534
rect 19997 14534 20080 14548
rect 19997 14522 20010 14534
rect 19568 14494 20010 14522
rect 19568 14482 19579 14494
rect 19505 14471 19579 14482
rect 19997 14482 20010 14494
rect 20062 14482 20080 14534
rect 19997 14468 20080 14482
rect 19819 14428 19901 14441
rect 19819 14372 19832 14428
rect 19888 14372 19901 14428
rect 19819 14359 19901 14372
rect 19188 14208 19258 14222
rect 19188 14156 19196 14208
rect 19248 14196 19258 14208
rect 19823 14208 19897 14219
rect 19823 14196 19834 14208
rect 19248 14168 19834 14196
rect 19248 14156 19258 14168
rect 13955 14138 14029 14149
rect 19188 14142 19258 14156
rect 19823 14156 19834 14168
rect 19886 14156 19897 14208
rect 19823 14145 19897 14156
rect 13955 14086 13966 14138
rect 14018 14086 14029 14138
rect 13955 14075 14029 14086
rect 13978 13739 14006 14075
rect 19765 14052 19847 14065
rect 19765 13996 19778 14052
rect 19834 13996 19847 14052
rect 19765 13983 19847 13996
rect 18146 13947 18382 13960
rect 13955 13728 14029 13739
rect 18146 13734 18154 13947
rect 18367 13937 20672 13947
rect 18367 13927 20675 13937
rect 18367 13734 20474 13927
rect 12914 13674 13478 13684
rect 13955 13676 13966 13728
rect 14018 13676 14029 13728
rect 20474 13716 20675 13726
rect 13955 13665 14029 13676
rect 19195 13636 19269 13647
rect 13858 13612 14096 13624
rect 13858 13560 13870 13612
rect 13922 13560 14030 13612
rect 14082 13560 14096 13612
rect 13858 13546 14096 13560
rect 14431 13614 14513 13627
rect 14431 13558 14444 13614
rect 14500 13558 14513 13614
rect 12914 13434 13478 13444
rect 13447 13312 13521 13323
rect 13447 13260 13458 13312
rect 13510 13260 13521 13312
rect 13447 13249 13521 13260
rect 12816 12470 13154 12492
rect 12816 12230 12840 12470
rect 13080 12230 13154 12470
rect 12816 12194 13154 12230
rect 13470 12169 13498 13249
rect 13950 13121 13978 13546
rect 14431 13545 14513 13558
rect 16287 13614 16369 13627
rect 16287 13558 16300 13614
rect 16356 13600 16369 13614
rect 16481 13612 16555 13623
rect 16481 13600 16492 13612
rect 16356 13572 16492 13600
rect 16356 13558 16369 13572
rect 16287 13545 16369 13558
rect 16481 13560 16492 13572
rect 16544 13560 16555 13612
rect 19195 13584 19206 13636
rect 19258 13584 19269 13636
rect 19195 13573 19269 13584
rect 16481 13549 16555 13560
rect 18391 13556 18465 13567
rect 18391 13544 18402 13556
rect 15361 13530 15435 13541
rect 15361 13478 15372 13530
rect 15424 13518 15435 13530
rect 15899 13530 15973 13541
rect 15899 13518 15910 13530
rect 15424 13490 15910 13518
rect 15424 13478 15435 13490
rect 15361 13467 15435 13478
rect 15899 13478 15910 13490
rect 15962 13478 15973 13530
rect 15899 13467 15973 13478
rect 18186 13516 18402 13544
rect 15278 13364 15356 13372
rect 15278 13312 15290 13364
rect 15342 13312 15356 13364
rect 15278 13306 15356 13312
rect 13927 13110 14001 13121
rect 13927 13058 13938 13110
rect 13990 13058 14001 13110
rect 13927 13047 14001 13058
rect 15302 13038 15330 13306
rect 18186 13151 18214 13516
rect 18391 13504 18402 13516
rect 18454 13504 18465 13556
rect 18391 13493 18465 13504
rect 19083 13476 19165 13489
rect 19218 13486 19246 13573
rect 19083 13420 19096 13476
rect 19152 13420 19165 13476
rect 19083 13407 19165 13420
rect 19194 13474 19270 13486
rect 19194 13422 19206 13474
rect 19258 13422 19270 13474
rect 19194 13410 19270 13422
rect 19101 13364 19175 13375
rect 19101 13312 19112 13364
rect 19164 13352 19175 13364
rect 19405 13364 19479 13375
rect 19405 13352 19416 13364
rect 19164 13324 19416 13352
rect 19164 13312 19175 13324
rect 19101 13301 19175 13312
rect 19405 13312 19416 13324
rect 19468 13312 19479 13364
rect 19405 13301 19479 13312
rect 19345 13232 19427 13245
rect 19047 13200 19129 13213
rect 18163 13140 18237 13151
rect 18163 13088 18174 13140
rect 18226 13088 18237 13140
rect 19047 13144 19060 13200
rect 19116 13144 19129 13200
rect 19345 13176 19358 13232
rect 19414 13176 19427 13232
rect 19345 13164 19427 13176
rect 19345 13163 19360 13164
rect 19047 13131 19129 13144
rect 19349 13112 19360 13163
rect 19412 13163 19427 13164
rect 19412 13112 19423 13163
rect 19349 13101 19423 13112
rect 18163 13077 18237 13088
rect 18857 13084 18931 13095
rect 15282 13032 15350 13038
rect 15282 12980 15290 13032
rect 15342 12980 15350 13032
rect 18857 13032 18868 13084
rect 18920 13072 18931 13084
rect 19056 13084 19120 13094
rect 19056 13072 19062 13084
rect 18920 13044 19062 13072
rect 18920 13032 18931 13044
rect 18857 13021 18931 13032
rect 19056 13032 19062 13044
rect 19114 13032 19120 13084
rect 19056 13022 19120 13032
rect 15282 12974 15350 12980
rect 18857 12978 18931 12989
rect 18857 12926 18868 12978
rect 18920 12966 18931 12978
rect 19071 12978 19145 12989
rect 19071 12966 19082 12978
rect 18920 12938 19082 12966
rect 18920 12926 18931 12938
rect 18857 12915 18931 12926
rect 19071 12926 19082 12938
rect 19134 12926 19145 12978
rect 19071 12915 19145 12926
rect 19349 12976 19423 12987
rect 19349 12924 19360 12976
rect 19412 12964 19423 12976
rect 19843 12976 19917 12987
rect 19843 12964 19854 12976
rect 19412 12936 19854 12964
rect 19412 12924 19423 12936
rect 19349 12913 19423 12924
rect 19843 12924 19854 12936
rect 19906 12924 19917 12976
rect 19843 12913 19917 12924
rect 21920 12913 22145 21553
rect 22416 21545 22425 21775
rect 22655 21545 22664 21775
rect 22978 21545 22987 21775
rect 23217 21545 23226 21775
rect 24066 21545 24075 21775
rect 24305 21545 24316 21775
rect 24626 21545 24635 21775
rect 24865 21545 24874 21775
rect 20208 12904 20416 12913
rect 15361 12866 15435 12877
rect 15361 12814 15372 12866
rect 15424 12854 15435 12866
rect 15424 12826 15978 12854
rect 15424 12814 15435 12826
rect 15361 12803 15435 12814
rect 13923 12768 14005 12783
rect 13923 12716 13938 12768
rect 13990 12716 14005 12768
rect 15950 12755 15978 12826
rect 16259 12824 16333 12835
rect 16259 12772 16270 12824
rect 16322 12812 16333 12824
rect 17179 12824 17253 12835
rect 17179 12812 17190 12824
rect 16322 12784 17190 12812
rect 16322 12772 16333 12784
rect 16259 12761 16333 12772
rect 17179 12772 17190 12784
rect 17242 12772 17253 12824
rect 17179 12761 17253 12772
rect 13923 12701 14005 12716
rect 15927 12744 16001 12755
rect 13447 12158 13521 12169
rect 13447 12106 13458 12158
rect 13510 12106 13521 12158
rect 13447 12095 13521 12106
rect 13950 11437 13978 12701
rect 15927 12692 15938 12744
rect 15990 12692 16001 12744
rect 18964 12740 18970 12861
rect 19091 12740 20208 12861
rect 15927 12681 16001 12692
rect 20208 12687 20416 12696
rect 21920 12679 22145 12688
rect 14624 12000 14718 12082
rect 17205 12080 17279 12089
rect 17205 12024 17210 12080
rect 17266 12078 17279 12080
rect 17268 12026 17279 12078
rect 17266 12024 17279 12026
rect 17205 12015 17279 12024
rect 19910 12082 20178 12100
rect 14624 11944 14638 12000
rect 14694 11944 14718 12000
rect 14624 11930 14718 11944
rect 17228 11677 17256 12015
rect 19349 11990 19423 12001
rect 17287 11974 17361 11985
rect 17287 11922 17298 11974
rect 17350 11962 17361 11974
rect 17795 11974 17869 11985
rect 17795 11962 17806 11974
rect 17350 11934 17806 11962
rect 17350 11922 17361 11934
rect 17287 11911 17361 11922
rect 17795 11922 17806 11934
rect 17858 11922 17869 11974
rect 19349 11938 19360 11990
rect 19412 11978 19423 11990
rect 19509 11990 19583 12001
rect 19509 11978 19520 11990
rect 19412 11950 19520 11978
rect 19412 11938 19423 11950
rect 19349 11927 19423 11938
rect 19509 11938 19520 11950
rect 19572 11938 19583 11990
rect 19509 11927 19583 11938
rect 17795 11911 17869 11922
rect 19910 11842 19922 12082
rect 20162 11842 20178 12082
rect 19910 11820 20178 11842
rect 17205 11666 17279 11677
rect 17205 11614 17216 11666
rect 17268 11614 17279 11666
rect 17205 11603 17279 11614
rect 13927 11426 14001 11437
rect 13927 11374 13938 11426
rect 13990 11374 14001 11426
rect 13927 11363 14001 11374
rect 16419 11174 16493 11185
rect 16419 11122 16430 11174
rect 16482 11122 16493 11174
rect 16419 11111 16493 11122
rect 16442 11025 16470 11111
rect 16789 11094 16863 11105
rect 16789 11042 16800 11094
rect 16852 11082 16863 11094
rect 17217 11094 17291 11105
rect 17217 11082 17228 11094
rect 16852 11054 17228 11082
rect 16852 11042 16863 11054
rect 16789 11031 16863 11042
rect 17217 11042 17228 11054
rect 17280 11042 17291 11094
rect 17217 11031 17291 11042
rect 16419 11014 16493 11025
rect 14567 10994 14641 11005
rect 13444 10942 13450 10994
rect 13502 10982 13508 10994
rect 14567 10982 14578 10994
rect 13502 10954 14578 10982
rect 13502 10942 13508 10954
rect 14567 10942 14578 10954
rect 14630 10942 14641 10994
rect 16419 10962 16430 11014
rect 16482 10962 16493 11014
rect 16419 10951 16493 10962
rect 14567 10931 14641 10942
rect 12774 10766 13044 10780
rect 12774 10526 12780 10766
rect 13020 10526 13044 10766
rect 12774 10510 13044 10526
rect 13593 10438 13667 10449
rect 13593 10386 13604 10438
rect 13656 10386 13667 10438
rect 13593 10375 13667 10386
rect 13616 9362 13644 10375
rect 14460 10242 14730 10260
rect 14460 10002 14476 10242
rect 14716 10002 14730 10242
rect 14460 9980 14730 10002
rect 19068 9470 19334 9480
rect 13837 9370 13911 9381
rect 13616 9334 13672 9362
rect 13369 9294 13443 9305
rect 13369 9242 13380 9294
rect 13432 9282 13443 9294
rect 13541 9294 13615 9305
rect 13541 9282 13552 9294
rect 13432 9254 13552 9282
rect 13432 9242 13443 9254
rect 13369 9231 13443 9242
rect 13541 9242 13552 9254
rect 13604 9242 13615 9294
rect 13541 9231 13615 9242
rect 13541 8306 13615 8317
rect 13288 8254 13294 8306
rect 13346 8294 13352 8306
rect 13541 8294 13552 8306
rect 13346 8266 13552 8294
rect 13346 8254 13352 8266
rect 13541 8254 13552 8266
rect 13604 8254 13615 8306
rect 13541 8243 13615 8254
rect 13369 8198 13443 8209
rect 13644 8198 13672 9334
rect 13837 9318 13848 9370
rect 13900 9318 13911 9370
rect 13837 9307 13911 9318
rect 13860 8209 13888 9307
rect 19068 8906 19334 8916
rect 14049 8304 14123 8315
rect 14049 8252 14060 8304
rect 14112 8292 14123 8304
rect 14273 8304 14347 8315
rect 14273 8292 14284 8304
rect 14112 8264 14284 8292
rect 14112 8252 14123 8264
rect 14049 8241 14123 8252
rect 14273 8252 14284 8264
rect 14336 8252 14347 8304
rect 14273 8241 14347 8252
rect 13369 8146 13380 8198
rect 13432 8186 13443 8198
rect 13594 8186 13600 8198
rect 13432 8158 13600 8186
rect 13432 8146 13443 8158
rect 13594 8146 13600 8158
rect 13652 8146 13672 8198
rect 13837 8198 13911 8209
rect 13837 8146 13848 8198
rect 13900 8146 13911 8198
rect 13369 8135 13443 8146
rect 13837 8135 13911 8146
rect 13627 7980 13709 7993
rect 13627 7924 13640 7980
rect 13696 7924 13709 7980
rect 13627 7911 13709 7924
rect 13860 7650 13888 8135
rect 14083 7980 14165 7993
rect 14083 7924 14096 7980
rect 14152 7924 14165 7980
rect 14083 7911 14165 7924
rect 13972 7650 13978 7662
rect 13860 7622 13978 7650
rect 13972 7610 13978 7622
rect 14030 7610 14036 7662
rect 14841 7160 14915 7171
rect 14841 7108 14852 7160
rect 14904 7148 14915 7160
rect 15033 7160 15107 7171
rect 15033 7148 15044 7160
rect 14904 7120 15044 7148
rect 14904 7108 14915 7120
rect 14841 7097 14915 7108
rect 15033 7108 15044 7120
rect 15096 7108 15107 7160
rect 15033 7097 15107 7108
rect 15927 7160 16001 7171
rect 15927 7108 15938 7160
rect 15990 7148 16001 7160
rect 16089 7160 16163 7171
rect 16089 7148 16100 7160
rect 15990 7120 16100 7148
rect 15990 7108 16001 7120
rect 15927 7097 16001 7108
rect 16089 7108 16100 7120
rect 16152 7108 16163 7160
rect 16089 7097 16163 7108
rect 17027 6764 17101 6775
rect 17027 6712 17038 6764
rect 17090 6712 17101 6764
rect 17027 6701 17101 6712
rect 17050 6455 17078 6701
rect 17027 6444 17101 6455
rect 17027 6392 17038 6444
rect 17090 6392 17101 6444
rect 17027 6381 17101 6392
rect 18153 6360 18227 6371
rect 18153 6308 18164 6360
rect 18216 6308 18227 6360
rect 18153 6297 18227 6308
rect 13060 5848 14898 5858
rect 17281 5528 17355 5539
rect 17281 5476 17292 5528
rect 17344 5476 17355 5528
rect 17281 5465 17355 5476
rect 13060 5424 14898 5434
rect 16251 5144 16325 5155
rect 16251 5092 16262 5144
rect 16314 5132 16325 5144
rect 17169 5144 17243 5155
rect 17169 5132 17180 5144
rect 16314 5104 17180 5132
rect 16314 5092 16325 5104
rect 16251 5081 16325 5092
rect 17169 5092 17180 5104
rect 17232 5092 17243 5144
rect 17169 5081 17243 5092
rect 17304 4839 17332 5465
rect 18176 5275 18204 6297
rect 18153 5264 18227 5275
rect 18153 5212 18164 5264
rect 18216 5212 18227 5264
rect 18153 5201 18227 5212
rect 17281 4828 17355 4839
rect 17281 4776 17292 4828
rect 17344 4776 17355 4828
rect 17281 4765 17355 4776
rect 18176 4664 18204 5201
rect 18152 4658 18228 4664
rect 18152 4606 18164 4658
rect 18216 4606 18228 4658
rect 13840 4584 13892 4590
rect 15575 4584 15649 4595
rect 18152 4594 18228 4606
rect 14978 4572 14984 4584
rect 13892 4544 14984 4572
rect 14978 4532 14984 4544
rect 15036 4572 15042 4584
rect 15575 4572 15586 4584
rect 15036 4544 15586 4572
rect 15036 4532 15042 4544
rect 15575 4532 15586 4544
rect 15638 4532 15649 4584
rect 13840 4526 13892 4532
rect 15575 4521 15649 4532
rect 14759 4376 14841 4391
rect 14759 4324 14774 4376
rect 14826 4324 14841 4376
rect 14759 4309 14841 4324
rect 13707 3634 13781 3645
rect 13707 3582 13718 3634
rect 13770 3582 13781 3634
rect 13707 3571 13781 3582
rect 13730 2771 13758 3571
rect 14786 3311 14814 4309
rect 17361 3986 17435 3997
rect 17361 3934 17372 3986
rect 17424 3934 17435 3986
rect 17361 3923 17435 3934
rect 17384 3649 17412 3923
rect 18176 3667 18204 4594
rect 19046 3698 19726 3708
rect 18153 3656 18227 3667
rect 17361 3638 17435 3649
rect 17361 3586 17372 3638
rect 17424 3586 17435 3638
rect 18153 3604 18164 3656
rect 18216 3604 18227 3656
rect 18153 3593 18227 3604
rect 17361 3575 17435 3586
rect 17366 3324 17372 3376
rect 17424 3324 17430 3376
rect 14763 3300 14837 3311
rect 14763 3248 14774 3300
rect 14826 3248 14837 3300
rect 14763 3237 14837 3248
rect 15075 3140 15149 3151
rect 15075 3088 15086 3140
rect 15138 3088 15149 3140
rect 15075 3077 15149 3088
rect 13707 2760 13781 2771
rect 13707 2708 13718 2760
rect 13770 2708 13781 2760
rect 13707 2697 13781 2708
rect 15098 2693 15126 3077
rect 15992 2848 16168 2858
rect 13819 2680 13893 2691
rect 13819 2628 13830 2680
rect 13882 2628 13893 2680
rect 13819 2617 13893 2628
rect 15075 2682 15149 2693
rect 15075 2630 15086 2682
rect 15138 2630 15149 2682
rect 15075 2619 15149 2630
rect 13707 2520 13781 2531
rect 13707 2468 13718 2520
rect 13770 2468 13781 2520
rect 13707 2457 13781 2468
rect 13730 1949 13758 2457
rect 13842 2283 13870 2617
rect 14897 2600 14971 2611
rect 14897 2548 14908 2600
rect 14960 2588 14971 2600
rect 15183 2600 15257 2611
rect 15183 2588 15194 2600
rect 14960 2560 15194 2588
rect 14960 2548 14971 2560
rect 14897 2537 14971 2548
rect 15183 2548 15194 2560
rect 15246 2548 15257 2600
rect 15183 2537 15257 2548
rect 15992 2378 16168 2388
rect 17384 2293 17412 3324
rect 19046 2958 19726 2968
rect 13819 2272 13893 2283
rect 13819 2220 13830 2272
rect 13882 2220 13893 2272
rect 13819 2209 13893 2220
rect 17357 2278 17439 2293
rect 17357 2226 17372 2278
rect 17424 2226 17439 2278
rect 17357 2211 17439 2226
rect 16251 2120 16325 2131
rect 16251 2068 16262 2120
rect 16314 2108 16325 2120
rect 16413 2120 16487 2131
rect 16413 2108 16424 2120
rect 16314 2080 16424 2108
rect 16314 2068 16325 2080
rect 16251 2057 16325 2068
rect 16413 2068 16424 2080
rect 16476 2068 16487 2120
rect 16413 2057 16487 2068
rect 13707 1938 13781 1949
rect 13707 1886 13718 1938
rect 13770 1886 13781 1938
rect 13707 1875 13781 1886
rect 18290 1780 18562 1800
rect 22420 1780 22660 21545
rect 22978 10280 23222 21545
rect 24070 16680 24316 21545
rect 24060 16665 24328 16680
rect 24060 16435 24081 16665
rect 24311 16435 24328 16665
rect 24060 16420 24328 16435
rect 24081 15156 24311 15160
rect 24076 15151 24316 15156
rect 24076 14921 24081 15151
rect 24311 14921 24316 15151
rect 22978 10239 23221 10280
rect 22978 10006 22983 10239
rect 23216 10006 23221 10239
rect 22978 10001 23221 10006
rect 22983 9997 23216 10001
rect 18290 1540 18306 1780
rect 18546 1540 18562 1780
rect 22411 1540 22420 1780
rect 22660 1540 22669 1780
rect 24076 1766 24316 14921
rect 24630 12470 24870 21545
rect 25162 21541 25171 21779
rect 25409 21541 25418 21779
rect 25166 13980 25414 21541
rect 25698 21538 25707 21782
rect 25951 21538 25960 21782
rect 25166 13723 25414 13732
rect 24630 12221 24870 12230
rect 25702 10793 25956 21538
rect 25702 10530 25956 10539
rect 18290 1514 18562 1540
rect 24076 1517 24316 1526
<< via2 >>
rect 4550 22150 4610 22210
rect 5092 22193 5148 22249
rect 5632 22192 5688 22248
rect 6212 22192 6268 22248
rect 6752 22192 6808 22248
rect 7332 22192 7388 22248
rect 7872 22192 7928 22248
rect 8432 22192 8488 22248
rect 8992 22192 9048 22248
rect 9552 22192 9608 22248
rect 10132 22192 10188 22248
rect 10672 22192 10728 22248
rect 11192 22192 11248 22248
rect 11752 22192 11808 22248
rect 12312 22192 12368 22248
rect 12872 22192 12928 22248
rect 13412 22192 13468 22248
rect 13972 22192 14028 22248
rect 14552 22192 14608 22248
rect 15072 22192 15128 22248
rect 15632 22192 15688 22248
rect 16172 22192 16228 22248
rect 16712 22192 16768 22248
rect 17272 22192 17328 22248
rect 21925 21553 22140 21768
rect 18992 16846 20700 20722
rect 19860 16450 20050 16650
rect 19358 15522 19414 15524
rect 19358 15470 19360 15522
rect 19360 15470 19412 15522
rect 19412 15470 19414 15522
rect 19358 15468 19414 15470
rect 19832 14426 19888 14428
rect 19832 14374 19834 14426
rect 19834 14374 19886 14426
rect 19886 14374 19888 14426
rect 19832 14372 19888 14374
rect 19778 14048 19834 14052
rect 19778 13996 19780 14048
rect 19780 13996 19832 14048
rect 19832 13996 19834 14048
rect 20474 13854 20675 13927
rect 20474 13802 20546 13854
rect 20546 13802 20598 13854
rect 20598 13802 20675 13854
rect 12914 13444 13478 13674
rect 20474 13726 20675 13802
rect 14444 13612 14500 13614
rect 14444 13560 14446 13612
rect 14446 13560 14498 13612
rect 14498 13560 14500 13612
rect 14444 13558 14500 13560
rect 12845 12235 13075 12465
rect 16300 13558 16356 13614
rect 19096 13474 19152 13476
rect 19096 13422 19098 13474
rect 19098 13422 19150 13474
rect 19150 13422 19152 13474
rect 19096 13420 19152 13422
rect 19060 13198 19116 13200
rect 19060 13146 19062 13198
rect 19062 13146 19114 13198
rect 19114 13146 19116 13198
rect 19060 13144 19116 13146
rect 19358 13176 19414 13232
rect 22425 21545 22655 21775
rect 22987 21545 23217 21775
rect 24075 21545 24305 21775
rect 24635 21545 24865 21775
rect 20208 12696 20416 12904
rect 21920 12688 22145 12913
rect 17210 12078 17266 12080
rect 17210 12026 17216 12078
rect 17216 12026 17266 12078
rect 17210 12024 17266 12026
rect 14638 11998 14694 12000
rect 14638 11946 14640 11998
rect 14640 11946 14692 11998
rect 14692 11946 14694 11998
rect 14638 11944 14694 11946
rect 19927 11847 20157 12077
rect 12785 10531 13015 10761
rect 14481 10007 14711 10237
rect 19068 8916 19334 9470
rect 13640 7978 13696 7980
rect 13640 7926 13642 7978
rect 13642 7926 13694 7978
rect 13694 7926 13696 7978
rect 13640 7924 13696 7926
rect 14096 7978 14152 7980
rect 14096 7926 14098 7978
rect 14098 7926 14150 7978
rect 14150 7926 14152 7978
rect 14096 7924 14152 7926
rect 13060 5434 14898 5848
rect 15992 2388 16168 2848
rect 19046 2968 19726 3698
rect 24081 16435 24311 16665
rect 24081 14921 24311 15151
rect 22983 10006 23216 10239
rect 18311 1545 18541 1775
rect 22420 1540 22660 1780
rect 25171 21541 25409 21779
rect 25707 21538 25951 21782
rect 25166 13732 25414 13980
rect 24630 12230 24870 12470
rect 25702 10539 25956 10793
rect 24076 1526 24316 1766
<< metal3 >>
rect 22956 22302 23236 22304
rect 21890 22298 22170 22300
rect 5060 22253 5180 22280
rect 4520 22214 4640 22240
rect 4520 22146 4546 22214
rect 4614 22146 4640 22214
rect 5060 22189 5088 22253
rect 5152 22189 5180 22253
rect 5060 22160 5180 22189
rect 5600 22252 5720 22280
rect 5600 22188 5628 22252
rect 5692 22188 5720 22252
rect 5600 22160 5720 22188
rect 6180 22252 6300 22280
rect 6180 22188 6208 22252
rect 6272 22188 6300 22252
rect 6180 22160 6300 22188
rect 6720 22252 6840 22280
rect 6720 22188 6748 22252
rect 6812 22188 6840 22252
rect 6720 22160 6840 22188
rect 7300 22252 7420 22280
rect 7300 22188 7328 22252
rect 7392 22188 7420 22252
rect 7300 22160 7420 22188
rect 7840 22252 7960 22280
rect 7840 22188 7868 22252
rect 7932 22188 7960 22252
rect 7840 22160 7960 22188
rect 8400 22252 8520 22280
rect 8400 22188 8428 22252
rect 8492 22188 8520 22252
rect 8400 22160 8520 22188
rect 8960 22252 9080 22280
rect 8960 22188 8988 22252
rect 9052 22188 9080 22252
rect 8960 22160 9080 22188
rect 9520 22252 9640 22280
rect 9520 22188 9548 22252
rect 9612 22188 9640 22252
rect 9520 22160 9640 22188
rect 10100 22252 10220 22280
rect 10100 22188 10128 22252
rect 10192 22188 10220 22252
rect 10100 22160 10220 22188
rect 10640 22252 10760 22280
rect 10640 22188 10668 22252
rect 10732 22188 10760 22252
rect 10640 22160 10760 22188
rect 11160 22252 11280 22280
rect 11160 22188 11188 22252
rect 11252 22188 11280 22252
rect 11160 22160 11280 22188
rect 11720 22252 11840 22280
rect 11720 22188 11748 22252
rect 11812 22188 11840 22252
rect 11720 22160 11840 22188
rect 12280 22252 12400 22280
rect 12280 22188 12308 22252
rect 12372 22188 12400 22252
rect 12280 22160 12400 22188
rect 12840 22252 12960 22280
rect 12840 22188 12868 22252
rect 12932 22188 12960 22252
rect 12840 22160 12960 22188
rect 13380 22252 13500 22280
rect 13380 22188 13408 22252
rect 13472 22188 13500 22252
rect 13380 22160 13500 22188
rect 13940 22252 14060 22280
rect 13940 22188 13968 22252
rect 14032 22188 14060 22252
rect 13940 22160 14060 22188
rect 14520 22252 14640 22280
rect 14520 22188 14548 22252
rect 14612 22188 14640 22252
rect 14520 22160 14640 22188
rect 15040 22252 15160 22280
rect 15040 22188 15068 22252
rect 15132 22188 15160 22252
rect 15040 22160 15160 22188
rect 15600 22252 15720 22280
rect 15600 22188 15628 22252
rect 15692 22188 15720 22252
rect 15600 22160 15720 22188
rect 16140 22252 16260 22280
rect 16140 22188 16168 22252
rect 16232 22188 16260 22252
rect 16140 22160 16260 22188
rect 16680 22252 16800 22280
rect 16680 22188 16708 22252
rect 16772 22188 16800 22252
rect 16680 22160 16800 22188
rect 17240 22252 17360 22280
rect 17240 22188 17268 22252
rect 17332 22188 17360 22252
rect 17240 22160 17360 22188
rect 4520 22120 4640 22146
rect 21890 22105 21939 22298
rect 22132 22105 22170 22298
rect 21890 22080 22170 22105
rect 22400 22280 22680 22300
rect 22400 22100 22420 22280
rect 22660 22100 22680 22280
rect 22956 22125 23011 22302
rect 23188 22125 23236 22302
rect 22956 22104 23236 22125
rect 24050 22296 24340 22300
rect 24050 22104 24104 22296
rect 24296 22104 24340 22296
rect 22400 22080 22680 22100
rect 21920 21770 22150 22080
rect 22420 21775 22660 22080
rect 21920 21768 22145 21770
rect 21920 21553 21925 21768
rect 22140 21553 22145 21768
rect 21920 21548 22145 21553
rect 22420 21545 22425 21775
rect 22655 21545 22660 21775
rect 22420 21540 22660 21545
rect 22982 21775 23222 22104
rect 24050 22100 24340 22104
rect 24608 22290 24894 22304
rect 25270 22300 25330 22304
rect 25686 22300 25968 22306
rect 24608 22100 24660 22290
rect 24830 22100 24894 22290
rect 22982 21545 22987 21775
rect 23217 21545 23222 21775
rect 22982 21540 23222 21545
rect 24070 21775 24310 22100
rect 24608 22088 24894 22100
rect 25150 22270 25430 22300
rect 25150 22100 25190 22270
rect 25390 22100 25430 22270
rect 25150 22090 25430 22100
rect 25686 22094 25720 22300
rect 25702 22092 25720 22094
rect 25942 22094 25968 22300
rect 25942 22092 25956 22094
rect 24070 21545 24075 21775
rect 24305 21545 24310 21775
rect 24070 21540 24310 21545
rect 24630 21775 24870 22088
rect 24630 21545 24635 21775
rect 24865 21545 24870 21775
rect 24630 21540 24870 21545
rect 25166 21779 25414 22090
rect 25166 21541 25171 21779
rect 25409 21541 25414 21779
rect 25166 21536 25414 21541
rect 25702 21782 25956 22092
rect 25702 21538 25707 21782
rect 25951 21538 25956 21782
rect 25702 21533 25956 21538
rect 18982 20722 20710 20727
rect 18982 16846 18992 20722
rect 20700 16846 20710 20722
rect 18982 16841 20710 16846
rect 24060 16670 24328 16680
rect 19836 16665 24328 16670
rect 19836 16650 24081 16665
rect 19836 16450 19860 16650
rect 20050 16450 24081 16650
rect 19836 16435 24081 16450
rect 24311 16435 24328 16665
rect 19836 16430 24328 16435
rect 24060 16420 24328 16430
rect 19346 15524 19427 15537
rect 19346 15468 19358 15524
rect 19414 15468 19427 15524
rect 19346 15455 19427 15468
rect 19356 15156 19416 15455
rect 19356 15151 24316 15156
rect 19356 14921 24081 15151
rect 24311 15121 24316 15151
rect 24311 14952 24318 15121
rect 24311 14921 24316 14952
rect 19356 14916 24316 14921
rect 12904 13674 13488 13679
rect 12904 13444 12914 13674
rect 13478 13444 13488 13674
rect 14431 13616 14513 13627
rect 16287 13616 16369 13627
rect 14431 13614 16369 13616
rect 14431 13558 14444 13614
rect 14500 13558 16300 13614
rect 16356 13558 16369 13614
rect 14431 13556 16369 13558
rect 14431 13545 14513 13556
rect 16287 13545 16369 13556
rect 12904 13439 13488 13444
rect 19083 13476 19165 13489
rect 19083 13420 19096 13476
rect 19152 13420 19165 13476
rect 19083 13407 19165 13420
rect 19094 13213 19154 13407
rect 19356 13245 19416 14916
rect 19819 14428 19901 14441
rect 19819 14372 19832 14428
rect 19888 14372 19901 14428
rect 19819 14359 19901 14372
rect 19830 14065 19890 14359
rect 19765 14052 19890 14065
rect 19765 13996 19778 14052
rect 19834 13996 19890 14052
rect 19765 13994 19890 13996
rect 19765 13983 19847 13994
rect 25161 13980 25419 13985
rect 20464 13929 20685 13932
rect 25161 13929 25166 13980
rect 20464 13927 25166 13929
rect 20464 13726 20474 13927
rect 20675 13732 25166 13927
rect 25414 13732 25419 13980
rect 20675 13728 25419 13732
rect 20675 13726 20685 13728
rect 25161 13727 25419 13728
rect 20464 13721 20685 13726
rect 19047 13200 19154 13213
rect 19047 13144 19060 13200
rect 19116 13144 19154 13200
rect 19345 13232 19427 13245
rect 19345 13176 19358 13232
rect 19414 13176 19427 13232
rect 19345 13163 19427 13176
rect 19047 13142 19154 13144
rect 19047 13131 19129 13142
rect 21915 12913 22150 12918
rect 21915 12909 21920 12913
rect 20203 12904 21920 12909
rect 20203 12696 20208 12904
rect 20416 12696 21920 12904
rect 20203 12691 21920 12696
rect 21915 12688 21920 12691
rect 22145 12909 22150 12913
rect 22145 12691 22160 12909
rect 22145 12688 22150 12691
rect 21915 12683 22150 12688
rect 12816 12470 13154 12492
rect 24625 12470 24875 12475
rect 12816 12465 24630 12470
rect 12816 12235 12845 12465
rect 13075 12235 24630 12465
rect 12816 12230 24630 12235
rect 24870 12230 24875 12470
rect 12816 12194 13154 12230
rect 24625 12225 24875 12230
rect 17205 12082 17271 12085
rect 14624 12080 17271 12082
rect 14624 12024 17210 12080
rect 17266 12024 17271 12080
rect 14624 12022 17271 12024
rect 14624 12000 14718 12022
rect 17205 12019 17271 12022
rect 19910 12082 20178 12100
rect 19910 12077 21512 12082
rect 14624 11944 14638 12000
rect 14694 11944 14718 12000
rect 14624 11930 14718 11944
rect 19910 11847 19927 12077
rect 20157 12073 21512 12077
rect 27550 12073 27781 12078
rect 20157 11852 30584 12073
rect 20157 11847 21512 11852
rect 27550 11847 27781 11852
rect 30304 11847 30584 11852
rect 19910 11842 21512 11847
rect 19910 11820 20178 11842
rect 25697 10793 25961 10798
rect 12774 10766 13044 10780
rect 12774 10761 21512 10766
rect 12774 10531 12785 10761
rect 13015 10753 21512 10761
rect 25697 10753 25702 10793
rect 13015 10539 25702 10753
rect 25956 10753 25961 10793
rect 25956 10539 25962 10753
rect 13015 10531 21512 10539
rect 25697 10534 25961 10539
rect 12774 10526 21512 10531
rect 12774 10510 13044 10526
rect 14460 10242 14730 10260
rect 15316 10242 23221 10244
rect 14460 10239 23221 10242
rect 14460 10237 22983 10239
rect 14460 10007 14481 10237
rect 14711 10007 22983 10237
rect 14460 10006 22983 10007
rect 23216 10006 23221 10239
rect 14460 10002 23221 10006
rect 14460 9980 14730 10002
rect 15316 10001 23221 10002
rect 19058 9470 19344 9475
rect 19058 8916 19068 9470
rect 19334 8916 19344 9470
rect 19058 8911 19344 8916
rect 13627 7982 13709 7993
rect 14083 7982 14165 7993
rect 13627 7980 14165 7982
rect 13627 7924 13640 7980
rect 13696 7924 14096 7980
rect 14152 7924 14165 7980
rect 13627 7922 14165 7924
rect 13627 7911 13709 7922
rect 14083 7911 14165 7922
rect 13050 5848 14908 5853
rect 13050 5434 13060 5848
rect 14898 5434 14908 5848
rect 13050 5429 14908 5434
rect 19036 3698 19736 3703
rect 19036 2968 19046 3698
rect 19726 2968 19736 3698
rect 19036 2963 19736 2968
rect 15982 2848 16178 2853
rect 15982 2388 15992 2848
rect 16168 2388 16178 2848
rect 15982 2383 16178 2388
rect 18290 1780 18562 1800
rect 22415 1780 22665 1785
rect 18290 1775 22420 1780
rect 18290 1545 18311 1775
rect 18541 1545 22420 1775
rect 18290 1540 22420 1545
rect 22660 1540 22665 1780
rect 18290 1514 18562 1540
rect 22415 1535 22665 1540
rect 24071 1766 24321 1771
rect 24071 1526 24076 1766
rect 24316 1750 25818 1766
rect 24316 1526 26372 1750
rect 24071 1521 24321 1526
rect 26098 190 26366 1526
rect 26098 70 26160 190
rect 26280 92 26366 190
rect 30306 200 30584 11847
rect 26280 70 26364 92
rect 26098 -2 26364 70
rect 30306 80 30392 200
rect 30512 80 30584 200
rect 30306 0 30584 80
<< via3 >>
rect 4546 22210 4614 22214
rect 4546 22150 4550 22210
rect 4550 22150 4610 22210
rect 4610 22150 4614 22210
rect 4546 22146 4614 22150
rect 5088 22249 5152 22253
rect 5088 22193 5092 22249
rect 5092 22193 5148 22249
rect 5148 22193 5152 22249
rect 5088 22189 5152 22193
rect 5628 22248 5692 22252
rect 5628 22192 5632 22248
rect 5632 22192 5688 22248
rect 5688 22192 5692 22248
rect 5628 22188 5692 22192
rect 6208 22248 6272 22252
rect 6208 22192 6212 22248
rect 6212 22192 6268 22248
rect 6268 22192 6272 22248
rect 6208 22188 6272 22192
rect 6748 22248 6812 22252
rect 6748 22192 6752 22248
rect 6752 22192 6808 22248
rect 6808 22192 6812 22248
rect 6748 22188 6812 22192
rect 7328 22248 7392 22252
rect 7328 22192 7332 22248
rect 7332 22192 7388 22248
rect 7388 22192 7392 22248
rect 7328 22188 7392 22192
rect 7868 22248 7932 22252
rect 7868 22192 7872 22248
rect 7872 22192 7928 22248
rect 7928 22192 7932 22248
rect 7868 22188 7932 22192
rect 8428 22248 8492 22252
rect 8428 22192 8432 22248
rect 8432 22192 8488 22248
rect 8488 22192 8492 22248
rect 8428 22188 8492 22192
rect 8988 22248 9052 22252
rect 8988 22192 8992 22248
rect 8992 22192 9048 22248
rect 9048 22192 9052 22248
rect 8988 22188 9052 22192
rect 9548 22248 9612 22252
rect 9548 22192 9552 22248
rect 9552 22192 9608 22248
rect 9608 22192 9612 22248
rect 9548 22188 9612 22192
rect 10128 22248 10192 22252
rect 10128 22192 10132 22248
rect 10132 22192 10188 22248
rect 10188 22192 10192 22248
rect 10128 22188 10192 22192
rect 10668 22248 10732 22252
rect 10668 22192 10672 22248
rect 10672 22192 10728 22248
rect 10728 22192 10732 22248
rect 10668 22188 10732 22192
rect 11188 22248 11252 22252
rect 11188 22192 11192 22248
rect 11192 22192 11248 22248
rect 11248 22192 11252 22248
rect 11188 22188 11252 22192
rect 11748 22248 11812 22252
rect 11748 22192 11752 22248
rect 11752 22192 11808 22248
rect 11808 22192 11812 22248
rect 11748 22188 11812 22192
rect 12308 22248 12372 22252
rect 12308 22192 12312 22248
rect 12312 22192 12368 22248
rect 12368 22192 12372 22248
rect 12308 22188 12372 22192
rect 12868 22248 12932 22252
rect 12868 22192 12872 22248
rect 12872 22192 12928 22248
rect 12928 22192 12932 22248
rect 12868 22188 12932 22192
rect 13408 22248 13472 22252
rect 13408 22192 13412 22248
rect 13412 22192 13468 22248
rect 13468 22192 13472 22248
rect 13408 22188 13472 22192
rect 13968 22248 14032 22252
rect 13968 22192 13972 22248
rect 13972 22192 14028 22248
rect 14028 22192 14032 22248
rect 13968 22188 14032 22192
rect 14548 22248 14612 22252
rect 14548 22192 14552 22248
rect 14552 22192 14608 22248
rect 14608 22192 14612 22248
rect 14548 22188 14612 22192
rect 15068 22248 15132 22252
rect 15068 22192 15072 22248
rect 15072 22192 15128 22248
rect 15128 22192 15132 22248
rect 15068 22188 15132 22192
rect 15628 22248 15692 22252
rect 15628 22192 15632 22248
rect 15632 22192 15688 22248
rect 15688 22192 15692 22248
rect 15628 22188 15692 22192
rect 16168 22248 16232 22252
rect 16168 22192 16172 22248
rect 16172 22192 16228 22248
rect 16228 22192 16232 22248
rect 16168 22188 16232 22192
rect 16708 22248 16772 22252
rect 16708 22192 16712 22248
rect 16712 22192 16768 22248
rect 16768 22192 16772 22248
rect 16708 22188 16772 22192
rect 17268 22248 17332 22252
rect 17268 22192 17272 22248
rect 17272 22192 17328 22248
rect 17328 22192 17332 22248
rect 17268 22188 17332 22192
rect 21939 22105 22132 22298
rect 22420 22100 22660 22280
rect 23011 22125 23188 22302
rect 24104 22104 24296 22296
rect 24660 22100 24830 22290
rect 25190 22100 25390 22270
rect 25720 22092 25942 22300
rect 18992 16846 20700 20722
rect 12914 13444 13478 13674
rect 19068 8916 19334 9470
rect 19046 2968 19726 3698
rect 15992 2388 16168 2848
rect 26160 70 26280 190
rect 30392 80 30512 200
<< metal4 >>
rect 4294 22215 4354 22304
rect 4846 22255 4906 22304
rect 4841 22253 5155 22255
rect 4294 22214 4615 22215
rect 4294 22146 4546 22214
rect 4614 22146 4615 22214
rect 4841 22189 5088 22253
rect 5152 22189 5155 22253
rect 4841 22185 5155 22189
rect 5398 22250 5458 22304
rect 5627 22252 5693 22253
rect 5627 22250 5628 22252
rect 5398 22190 5628 22250
rect 4294 22145 4615 22146
rect 4294 22104 4354 22145
rect 4846 22104 4906 22185
rect 5398 22104 5458 22190
rect 5627 22188 5628 22190
rect 5692 22188 5693 22252
rect 5627 22187 5693 22188
rect 5950 22250 6010 22304
rect 6207 22252 6273 22253
rect 6207 22250 6208 22252
rect 5950 22190 6208 22250
rect 5950 22104 6010 22190
rect 6207 22188 6208 22190
rect 6272 22188 6273 22252
rect 6207 22187 6273 22188
rect 6502 22250 6562 22304
rect 6747 22252 6813 22253
rect 6747 22250 6748 22252
rect 6502 22190 6748 22250
rect 6502 22104 6562 22190
rect 6747 22188 6748 22190
rect 6812 22188 6813 22252
rect 6747 22187 6813 22188
rect 7054 22250 7114 22304
rect 7327 22252 7393 22253
rect 7327 22250 7328 22252
rect 7054 22190 7328 22250
rect 7054 22104 7114 22190
rect 7327 22188 7328 22190
rect 7392 22188 7393 22252
rect 7327 22187 7393 22188
rect 7606 22250 7666 22304
rect 7867 22252 7933 22253
rect 7867 22250 7868 22252
rect 7606 22190 7868 22250
rect 7606 22104 7666 22190
rect 7867 22188 7868 22190
rect 7932 22188 7933 22252
rect 7867 22187 7933 22188
rect 8158 22250 8218 22304
rect 8427 22252 8493 22253
rect 8427 22250 8428 22252
rect 8158 22190 8428 22250
rect 8158 22104 8218 22190
rect 8427 22188 8428 22190
rect 8492 22188 8493 22252
rect 8427 22187 8493 22188
rect 8710 22250 8770 22304
rect 8987 22252 9053 22253
rect 8987 22250 8988 22252
rect 8710 22190 8988 22250
rect 8710 22104 8770 22190
rect 8987 22188 8988 22190
rect 9052 22188 9053 22252
rect 8987 22187 9053 22188
rect 9262 22250 9322 22304
rect 9547 22252 9613 22253
rect 9547 22250 9548 22252
rect 9262 22190 9548 22250
rect 9262 22104 9322 22190
rect 9547 22188 9548 22190
rect 9612 22188 9613 22252
rect 9547 22187 9613 22188
rect 9814 22250 9874 22304
rect 10127 22252 10193 22253
rect 10127 22250 10128 22252
rect 9814 22190 10128 22250
rect 9814 22104 9874 22190
rect 10127 22188 10128 22190
rect 10192 22188 10193 22252
rect 10127 22187 10193 22188
rect 10366 22250 10426 22304
rect 10667 22252 10733 22253
rect 10667 22250 10668 22252
rect 10366 22190 10668 22250
rect 10366 22104 10426 22190
rect 10667 22188 10668 22190
rect 10732 22188 10733 22252
rect 10667 22187 10733 22188
rect 10918 22250 10978 22304
rect 11187 22252 11253 22253
rect 11187 22250 11188 22252
rect 10918 22190 11188 22250
rect 10918 22104 10978 22190
rect 11187 22188 11188 22190
rect 11252 22188 11253 22252
rect 11187 22187 11253 22188
rect 11470 22250 11530 22304
rect 11747 22252 11813 22253
rect 11747 22250 11748 22252
rect 11470 22190 11748 22250
rect 11470 22104 11530 22190
rect 11747 22188 11748 22190
rect 11812 22188 11813 22252
rect 11747 22187 11813 22188
rect 12022 22250 12082 22304
rect 12307 22252 12373 22253
rect 12307 22250 12308 22252
rect 12022 22190 12308 22250
rect 12022 22104 12082 22190
rect 12307 22188 12308 22190
rect 12372 22188 12373 22252
rect 12307 22187 12373 22188
rect 12574 22250 12634 22304
rect 12867 22252 12933 22253
rect 12867 22250 12868 22252
rect 12574 22190 12868 22250
rect 12574 22104 12634 22190
rect 12867 22188 12868 22190
rect 12932 22188 12933 22252
rect 12867 22187 12933 22188
rect 13126 22250 13186 22304
rect 13407 22252 13473 22253
rect 13407 22250 13408 22252
rect 13126 22190 13408 22250
rect 13126 22104 13186 22190
rect 13407 22188 13408 22190
rect 13472 22188 13473 22252
rect 13407 22187 13473 22188
rect 13678 22250 13738 22304
rect 13967 22252 14033 22253
rect 13967 22250 13968 22252
rect 13678 22190 13968 22250
rect 13678 22104 13738 22190
rect 13967 22188 13968 22190
rect 14032 22188 14033 22252
rect 13967 22187 14033 22188
rect 14230 22250 14290 22304
rect 14547 22252 14613 22253
rect 14547 22250 14548 22252
rect 14230 22190 14548 22250
rect 14230 22104 14290 22190
rect 14547 22188 14548 22190
rect 14612 22188 14613 22252
rect 14547 22187 14613 22188
rect 14782 22250 14842 22304
rect 15067 22252 15133 22253
rect 15067 22250 15068 22252
rect 14782 22190 15068 22250
rect 14782 22104 14842 22190
rect 15067 22188 15068 22190
rect 15132 22188 15133 22252
rect 15067 22187 15133 22188
rect 15334 22250 15394 22304
rect 15627 22252 15693 22253
rect 15627 22250 15628 22252
rect 15334 22190 15628 22250
rect 15334 22104 15394 22190
rect 15627 22188 15628 22190
rect 15692 22188 15693 22252
rect 15627 22187 15693 22188
rect 15886 22250 15946 22304
rect 16167 22252 16233 22253
rect 16167 22250 16168 22252
rect 15886 22190 16168 22250
rect 15886 22104 15946 22190
rect 16167 22188 16168 22190
rect 16232 22188 16233 22252
rect 16167 22187 16233 22188
rect 16438 22250 16498 22304
rect 16707 22252 16773 22253
rect 16707 22250 16708 22252
rect 16438 22190 16708 22250
rect 16438 22104 16498 22190
rect 16707 22188 16708 22190
rect 16772 22188 16773 22252
rect 16707 22187 16773 22188
rect 16990 22250 17050 22304
rect 17267 22252 17333 22253
rect 17267 22250 17268 22252
rect 16990 22190 17268 22250
rect 16990 22104 17050 22190
rect 17267 22188 17268 22190
rect 17332 22188 17333 22252
rect 17267 22187 17333 22188
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 22299 22018 22304
rect 22510 22301 22570 22304
rect 23062 22303 23122 22304
rect 23010 22302 23189 22303
rect 21938 22298 22133 22299
rect 21938 22105 21939 22298
rect 22132 22105 22133 22298
rect 22500 22281 22580 22301
rect 21938 22104 22133 22105
rect 22419 22280 22661 22281
rect 22419 22100 22420 22280
rect 22660 22100 22661 22280
rect 23010 22125 23011 22302
rect 23188 22125 23189 22302
rect 23010 22124 23189 22125
rect 23010 22112 23188 22124
rect 23614 22104 23674 22304
rect 24166 22297 24226 22304
rect 24718 22298 24778 22304
rect 24103 22296 24297 22297
rect 24103 22104 24104 22296
rect 24296 22104 24297 22296
rect 24103 22103 24297 22104
rect 24652 22290 24840 22298
rect 22419 22099 22661 22100
rect 24652 22100 24660 22290
rect 24830 22100 24840 22290
rect 25270 22280 25330 22304
rect 25822 22301 25882 22304
rect 25719 22300 25943 22301
rect 24652 22094 24840 22100
rect 25180 22270 25400 22280
rect 25180 22100 25190 22270
rect 25390 22100 25400 22270
rect 25180 22090 25400 22100
rect 25719 22092 25720 22300
rect 25942 22092 25943 22300
rect 26374 22104 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 25719 22091 25943 22092
rect 11868 13674 17732 21658
rect 11868 13444 12914 13674
rect 13478 13444 17732 13674
rect 11868 2848 17732 13444
rect 11868 2388 15992 2848
rect 16168 2388 17732 2848
rect 11868 630 17732 2388
rect 18930 20722 24794 21604
rect 18930 16846 18992 20722
rect 20700 16846 24794 20722
rect 18930 9470 24794 16846
rect 18930 8916 19068 9470
rect 19334 8916 24794 9470
rect 18930 3698 24794 8916
rect 18930 2968 19046 3698
rect 19726 2968 24794 3698
rect 18930 576 24794 2968
rect 30391 200 30513 201
rect 768 0 888 200
rect 5000 0 5120 200
rect 9232 0 9352 200
rect 13464 0 13584 200
rect 17696 0 17816 200
rect 21928 0 22048 200
rect 26160 191 26280 200
rect 26159 190 26281 191
rect 26159 70 26160 190
rect 26280 70 26281 190
rect 30391 80 30392 200
rect 30512 80 30513 200
rect 30391 79 30513 80
rect 26159 69 26281 70
rect 26160 0 26280 69
rect 30392 0 30512 79
use XM1_xbuf1_xringosc  XM1_xbuf1_xringosc_0 dev
timestamp 1698067942
transform 0 1 14768 -1 0 2323
box -246 -1179 246 1179
use XM1_xbuf2_xringosc  XM1_xbuf2_xringosc_0 dev
timestamp 1698067942
transform 0 1 18207 -1 0 8729
box -246 -1179 246 1179
use XM1_xbuf3_xringosc  XM1_xbuf3_xringosc_0 dev
timestamp 1698067942
transform 0 1 15022 -1 0 7237
box -246 -1179 246 1179
use XM1_xdrv_b0_xdac  XM1_xdrv_b0_xdac_0 dev
timestamp 1698067942
transform 0 -1 13446 1 0 10987
box -246 -679 246 679
use XM1_xdrv_b1_xdac  XM1_xdrv_b1_xdac_0 dev
timestamp 1698067942
transform 0 1 17735 -1 0 13702
box -246 -679 246 679
use XM1_xdrv_b2_xdac  XM1_xdrv_b2_xdac_0 dev
timestamp 1698067942
transform -1 0 13976 0 -1 13171
box -246 -679 246 679
use XM1_xdrv_dummy_xdac  XM1_xdrv_dummy_xdac_0 dev
timestamp 1698067942
transform 0 1 17773 -1 0 11972
box -246 -679 246 679
use XM1_xro1_xringosc  XM1_xro1_xringosc_0 dev
timestamp 1698067942
transform -1 0 17397 0 -1 2173
box -1196 -234 1196 234
use XM1_xro2_xringosc  XM1_xro2_xringosc_0 dev
timestamp 1698067942
transform 1 0 18189 0 1 6419
box -1196 -234 1196 234
use XM1_xro3_xringosc  XM1_xro3_xringosc_0 dev
timestamp 1698067942
transform 0 -1 13824 1 0 4557
box -1196 -234 1196 234
use XM1_xtgbyp  XM1_xtgbyp_0 dev
timestamp 1698067942
transform 0 -1 19006 1 0 13357
box -246 -279 246 279
use XM1_xtgdac  XM1_xtgdac_0 dev
timestamp 1698067942
transform 0 1 19925 -1 0 14102
box -246 -279 246 279
use XM1_xtgro  XM1_xtgro_0 dev
timestamp 1698067942
transform 0 1 14198 -1 0 7872
box -246 -279 246 279
use XM2_xtgbyp  XM2_xtgbyp_0 dev
timestamp 1698067942
transform 0 -1 19670 1 0 13356
box -246 -384 246 384
use XM2_xtgdac  XM2_xtgdac_0 dev
timestamp 1698067942
transform 0 1 19261 -1 0 14103
box -246 -384 246 384
use XM2_xtgro  XM2_xtgro_0 dev
timestamp 1698067942
transform 0 1 13534 -1 0 7873
box -246 -384 246 384
use XM2A_xbuf1_xringosc  XM2A_xbuf1_xringosc_0 dev
timestamp 1698067942
transform 0 1 14762 -1 0 1831
box -246 -1184 246 1184
use XM2A_xbuf2_xringosc  XM2A_xbuf2_xringosc_0 dev
timestamp 1698067942
transform 0 1 18201 -1 0 8237
box -246 -1184 246 1184
use XM2A_xbuf3_xringosc  XM2A_xbuf3_xringosc_0 dev
timestamp 1698067942
transform 0 1 15016 -1 0 6745
box -246 -1184 246 1184
use XM2A_xdrv_b0_xdac  XM2A_xdrv_b0_xdac_0 dev
timestamp 1698067942
transform 0 -1 13430 1 0 11971
box -246 -684 246 684
use XM2A_xdrv_b1_xdac  XM2A_xdrv_b1_xdac_0 dev
timestamp 1698067942
transform 0 1 17751 -1 0 12718
box -246 -684 246 684
use XM2A_xdrv_b2_xdac  XM2A_xdrv_b2_xdac_0 dev
timestamp 1698067942
transform -1 0 12992 0 -1 13155
box -246 -684 246 684
use XM2A_xdrv_dummy_xdac  XM2A_xdrv_dummy_xdac_0 dev
timestamp 1698067942
transform 0 1 17789 -1 0 10988
box -246 -684 246 684
use XM2A_xro1_xringosc  XM2A_xro1_xringosc_0 dev
timestamp 1698067942
transform -1 0 17397 0 -1 3428
box -1196 -229 1196 229
use XM2A_xro2_xringosc  XM2A_xro2_xringosc_0 dev
timestamp 1698067942
transform 1 0 18189 0 1 5164
box -1196 -229 1196 229
use XM2A_xro3_xringosc  XM2A_xro3_xringosc_0 dev
timestamp 1698067942
transform 0 -1 15079 1 0 4557
box -1196 -229 1196 229
use XM2B_xbuf1_xringosc  XM2B_xbuf1_xringosc_0 dev
timestamp 1698067942
transform 0 1 14762 -1 0 1339
box -246 -1184 246 1184
use XM2B_xbuf2_xringosc  XM2B_xbuf2_xringosc_0 dev
timestamp 1698067942
transform 0 1 18201 -1 0 7745
box -246 -1184 246 1184
use XM2B_xbuf3_xringosc  XM2B_xbuf3_xringosc_0 dev
timestamp 1698067942
transform 0 1 15016 -1 0 6253
box -246 -1184 246 1184
use XM2B_xdrv_b0_xdac  XM2B_xdrv_b0_xdac_0 dev
timestamp 1698067942
transform 0 -1 13430 1 0 11479
box -246 -684 246 684
use XM2B_xdrv_b1_xdac  XM2B_xdrv_b1_xdac_0 dev
timestamp 1698067942
transform 0 1 17751 -1 0 13210
box -246 -684 246 684
use XM2B_xdrv_b2_xdac  XM2B_xdrv_b2_xdac_0 dev
timestamp 1698067942
transform -1 0 13484 0 -1 13155
box -246 -684 246 684
use XM2B_xdrv_dummy_xdac  XM2B_xdrv_dummy_xdac_0 dev
timestamp 1698067942
transform 0 1 17789 -1 0 11480
box -246 -684 246 684
use XM2B_xro1_xringosc  XM2B_xro1_xringosc_0 dev
timestamp 1698067942
transform 1 0 17397 0 1 3886
box -1196 -229 1196 229
use XM2B_xro2_xringosc  XM2B_xro2_xringosc_0 dev
timestamp 1698067942
transform -1 0 18189 0 -1 4706
box -1196 -229 1196 229
use XM2B_xro3_xringosc  XM2B_xro3_xringosc_0 dev
timestamp 1698067942
transform 0 1 15537 -1 0 4557
box -1196 -229 1196 229
use XM3_xdrv_b0_xdac  XM3_xdrv_b0_xdac_0 dev
timestamp 1698067942
transform 0 1 14804 -1 0 10987
box -246 -679 246 679
use XM3_xdrv_b1_xdac  XM3_xdrv_b1_xdac_0 dev
timestamp 1698067942
transform 0 -1 16377 1 0 13702
box -246 -679 246 679
use XM3_xdrv_b2_xdac  XM3_xdrv_b2_xdac_0 dev
timestamp 1698067942
transform 1 0 13976 0 1 14529
box -246 -679 246 679
use XM3_xdrv_dummy_xdac  XM3_xdrv_dummy_xdac_0 dev
timestamp 1698067942
transform 0 -1 16415 1 0 11972
box -246 -679 246 679
use XM3_xtgbyp  XM3_xtgbyp_0 dev
timestamp 1698067942
transform -1 0 18974 0 -1 11932
box -246 -1179 246 1179
use XM3_xtgdac  XM3_xtgdac_0 dev
timestamp 1698067942
transform 1 0 19957 0 1 15527
box -246 -1179 246 1179
use XM3_xtgro  XM3_xtgro_0 dev
timestamp 1698067942
transform 1 0 14230 0 1 9297
box -246 -1179 246 1179
use XM4A_xdrv_b0_xdac  XM4A_xdrv_b0_xdac_0 dev
timestamp 1698067942
transform 0 1 14798 -1 0 11479
box -246 -684 246 684
use XM4A_xdrv_b1_xdac  XM4A_xdrv_b1_xdac_0 dev
timestamp 1698067942
transform 0 -1 16383 1 0 13210
box -246 -684 246 684
use XM4A_xdrv_b2_xdac  XM4A_xdrv_b2_xdac_0 dev
timestamp 1698067942
transform 1 0 13484 0 1 14523
box -246 -684 246 684
use XM4A_xdrv_dummy_xdac  XM4A_xdrv_dummy_xdac_0 dev
timestamp 1698067942
transform 0 -1 16421 1 0 11480
box -246 -684 246 684
use XM4A_xtgbyp  XM4A_xtgbyp_0 dev
timestamp 1698067942
transform -1 0 19466 0 -1 11926
box -246 -1184 246 1184
use XM4A_xtgdac  XM4A_xtgdac_0 dev
timestamp 1698067942
transform 1 0 19465 0 1 15533
box -246 -1184 246 1184
use XM4A_xtgro  XM4A_xtgro_0 dev
timestamp 1698067942
transform 1 0 13738 0 1 9303
box -246 -1184 246 1184
use XM4B_xdrv_b0_xdac  XM4B_xdrv_b0_xdac_0 dev
timestamp 1698067942
transform 0 1 14798 -1 0 11971
box -246 -684 246 684
use XM4B_xdrv_b1_xdac  XM4B_xdrv_b1_xdac_0 dev
timestamp 1698067942
transform 0 -1 16383 1 0 12718
box -246 -684 246 684
use XM4B_xdrv_b2_xdac  XM4B_xdrv_b2_xdac_0 dev
timestamp 1698067942
transform 1 0 12992 0 1 14523
box -246 -684 246 684
use XM4B_xdrv_dummy_xdac  XM4B_xdrv_dummy_xdac_0 dev
timestamp 1698067942
transform 0 -1 16421 1 0 10988
box -246 -684 246 684
use XM4B_xtgbyp  XM4B_xtgbyp_0 dev
timestamp 1698067942
transform -1 0 19958 0 -1 11926
box -246 -1184 246 1184
use XM4B_xtgdac  XM4B_xtgdac_0 dev
timestamp 1698067942
transform 1 0 18973 0 1 15533
box -246 -1184 246 1184
use XM4B_xtgro  XM4B_xtgro_0 dev
timestamp 1698067942
transform 1 0 13246 0 1 9303
box -246 -1184 246 1184
use XMcap1_xro1_xringosc  XMcap1_xro1_xringosc_0 dev
timestamp 1698067942
transform -1 0 18989 0 -1 3117
box -396 -1179 396 1179
use XMcap1_xro2_xringosc  XMcap1_xro2_xringosc_0 dev
timestamp 1698067942
transform 1 0 16597 0 1 5475
box -396 -1179 396 1179
use XMcap1_xro3_xringosc  XMcap1_xro3_xringosc_0 dev
timestamp 1698067942
transform 0 -1 14768 1 0 2965
box -396 -1179 396 1179
use XMcap2_xro1_xringosc  XMcap2_xro1_xringosc_0 dev
timestamp 1698067942
transform 0 1 17385 -1 0 2803
box -396 -1184 396 1184
use XMcap2_xro2_xringosc  XMcap2_xro2_xringosc_0 dev
timestamp 1698067942
transform 0 -1 18201 1 0 5789
box -396 -1184 396 1184
use XMcap2_xro3_xringosc  XMcap2_xro3_xringosc_0 dev
timestamp 1698067942
transform -1 0 14454 0 -1 4569
box -396 -1184 396 1184
use XMpowerdn_xro1_xringosc  XMpowerdn_xro1_xringosc_0 dev
timestamp 1698067942
transform 0 1 17385 -1 0 1643
box -296 -1184 296 1184
use XMpowerdn_xro2_xringosc  XMpowerdn_xro2_xringosc_0 dev
timestamp 1698067942
transform 0 -1 18201 1 0 6949
box -296 -1184 296 1184
use XMpowerdn_xro3_xringosc  XMpowerdn_xro3_xringosc_0 dev
timestamp 1698067942
transform -1 0 13294 0 -1 4569
box -296 -1184 296 1184
use XR1  XR1_0 dev
timestamp 1698067942
transform 1 0 8461 0 1 21333
box -201 -633 201 633
use XR2  XR2_0 dev
timestamp 1698067942
transform 1 0 7901 0 1 21333
box -201 -633 201 633
use XR3  XR3_0 dev
timestamp 1698067942
transform 1 0 7361 0 1 21333
box -201 -633 201 633
use XR4  XR4_0 dev
timestamp 1698067942
transform 1 0 6781 0 1 21333
box -201 -633 201 633
use XR5  XR5_0 dev
timestamp 1698067942
transform 1 0 6241 0 1 21333
box -201 -633 201 633
use XR6  XR6_0 dev
timestamp 1698067942
transform 1 0 5661 0 1 21333
box -201 -633 201 633
use XR7  XR7_1 dev
timestamp 1698067942
transform 1 0 5121 0 1 21333
box -201 -633 201 633
use XR8  XR8_0 dev
timestamp 1698067942
transform 1 0 4581 0 1 21333
box -201 -633 201 633
use XR9  XR9_0 dev
timestamp 1698067942
transform 1 0 12901 0 1 21333
box -201 -633 201 633
use XR10  XR10_0 dev
timestamp 1698067942
transform 1 0 12341 0 1 21333
box -201 -633 201 633
use XR11  XR11_0 dev
timestamp 1698067942
transform 1 0 11781 0 1 21333
box -201 -633 201 633
use XR12  XR12_0 dev
timestamp 1698067942
transform 1 0 11221 0 1 21333
box -201 -633 201 633
use XR13  XR13_0 dev
timestamp 1698067942
transform 1 0 10701 0 1 21333
box -201 -633 201 633
use XR14  XR14_0 dev
timestamp 1698067942
transform 1 0 10161 0 1 21333
box -201 -633 201 633
use XR15  XR15_0 dev
timestamp 1698067942
transform 1 0 9581 0 1 21333
box -201 -633 201 633
use XR16  XR16_0 dev
timestamp 1698067942
transform 1 0 9021 0 1 21333
box -201 -633 201 633
use XR17  XR17_0 dev
timestamp 1698067942
transform 1 0 17301 0 1 21333
box -201 -633 201 633
use XR18  XR18_0 dev
timestamp 1698067942
transform 1 0 16741 0 1 21333
box -201 -633 201 633
use XR19  XR19_0 dev
timestamp 1698067942
transform 1 0 16201 0 1 21333
box -201 -633 201 633
use XR20  XR20_0 dev
timestamp 1698067942
transform 1 0 15661 0 1 21333
box -201 -633 201 633
use XR21  XR21_0 dev
timestamp 1698067942
transform 1 0 15101 0 1 21333
box -201 -633 201 633
use XR22  XR22_0 dev
timestamp 1698067942
transform 1 0 14581 0 1 21333
box -201 -633 201 633
use XR23  XR23_0 dev
timestamp 1698067942
transform 1 0 14001 0 1 21333
box -201 -633 201 633
use XR24  XR24_0 dev
timestamp 1698067942
transform 1 0 13441 0 1 21333
box -201 -633 201 633
use XRSTR_0_xdac  XRSTR_0_xdac_0 dev
timestamp 1698067942
transform 0 1 14960 -1 0 13586
box -1114 -738 1114 738
<< labels >>
flabel metal4 s 26926 22104 26986 22304 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 27478 22104 27538 22304 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 26374 22104 26434 22304 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30392 0 30512 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26160 0 26280 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 21928 0 22048 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 17696 0 17816 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13464 0 13584 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 5000 0 5120 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 768 0 888 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 24718 22104 24778 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 24166 22104 24226 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 23062 22104 23122 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21958 22104 22018 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 20854 22104 20914 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 20302 22104 20362 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 19750 22104 19810 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 18646 22104 18706 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 18094 22104 18154 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 17542 22104 17602 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 7606 22104 7666 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 7054 22104 7114 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 6502 22104 6562 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 5398 22104 5458 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 4846 22104 4906 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 4294 22104 4354 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 12022 22104 12082 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 11470 22104 11530 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 10918 22104 10978 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 9814 22104 9874 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 9262 22104 9322 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 8710 22104 8770 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16438 22104 16498 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 15886 22104 15946 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15334 22104 15394 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14230 22104 14290 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13678 22104 13738 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 13126 22104 13186 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 s 26926 22104 26986 22304 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 27478 22104 27538 22304 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 26374 22104 26434 22304 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30392 0 30512 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26160 0 26280 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 21928 0 22048 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 17696 0 17816 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13464 0 13584 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 5000 0 5120 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 768 0 888 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 25270 22104 25330 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 24718 22104 24778 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 24166 22104 24226 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 23062 22104 23122 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21958 22104 22018 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 20854 22104 20914 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 20302 22104 20362 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 19750 22104 19810 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 18646 22104 18706 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 18094 22104 18154 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 17542 22104 17602 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 7606 22104 7666 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 7054 22104 7114 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 6502 22104 6562 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 5398 22104 5458 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 4846 22104 4906 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 4294 22104 4354 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 12022 22104 12082 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 11470 22104 11530 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 10918 22104 10978 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 9814 22104 9874 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 9262 22104 9322 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 8710 22104 8770 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16438 22104 16498 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 15886 22104 15946 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15334 22104 15394 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14230 22104 14290 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13678 22104 13738 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 13126 22104 13186 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 s 22510 22104 22570 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 22510 22104 22570 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
rlabel metal4 11868 630 17732 21658 1 VPWR
rlabel metal4 18930 576 24794 21604 1 VGND
flabel metal4 14400 800 14800 21600 1 FreeSerif 3200 0 0 0 VPWR
port 51 n
flabel metal4 21600 800 22000 21600 1 FreeSerif 3200 0 0 0 VGND
port 52 n
<< properties >>
string FIXED_BBOX 0 0 31464 22304
<< end >>
