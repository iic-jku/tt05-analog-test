magic
tech sky130A
magscale 1 2
timestamp 1698067942
<< nwell >>
rect -396 -1184 396 1184
<< pmos >>
rect -200 -1036 200 964
<< pdiff >>
rect -258 952 -200 964
rect -258 -1024 -246 952
rect -212 -1024 -200 952
rect -258 -1036 -200 -1024
rect 200 952 258 964
rect 200 -1024 212 952
rect 246 -1024 258 952
rect 200 -1036 258 -1024
<< pdiffc >>
rect -246 -1024 -212 952
rect 212 -1024 246 952
<< nsubdiff >>
rect -360 1114 360 1148
rect -360 -1114 -326 1114
rect 326 -1114 360 1114
rect -360 -1148 -264 -1114
rect 264 -1148 360 -1114
<< nsubdiffcont >>
rect -264 -1148 264 -1114
<< poly >>
rect -200 1045 200 1061
rect -200 1011 -184 1045
rect 184 1011 200 1045
rect -200 964 200 1011
rect -200 -1062 200 -1036
<< polycont >>
rect -184 1011 184 1045
<< locali >>
rect -360 1114 360 1148
rect -360 -1114 -326 1114
rect -200 1011 -184 1045
rect 184 1011 200 1045
rect -246 952 -212 968
rect -246 -1040 -212 -1024
rect 212 952 246 968
rect 212 -1040 246 -1024
rect 326 -1114 360 1114
rect -360 -1148 -264 -1114
rect 264 -1148 360 -1114
<< properties >>
string FIXED_BBOX -343 -1131 343 1131
<< end >>
