magic
tech sky130A
magscale 1 2
timestamp 1698067942
<< nwell >>
rect -1196 -234 1196 234
<< pmos >>
rect -1000 -86 1000 14
<< pdiff >>
rect -1058 2 -1000 14
rect -1058 -74 -1046 2
rect -1012 -74 -1000 2
rect -1058 -86 -1000 -74
rect 1000 2 1058 14
rect 1000 -74 1012 2
rect 1046 -74 1058 2
rect 1000 -86 1058 -74
<< pdiffc >>
rect -1046 -74 -1012 2
rect 1012 -74 1046 2
<< nsubdiff >>
rect -1160 164 1160 198
rect -1160 -164 -1126 164
rect 1126 -164 1160 164
rect -1160 -198 -1064 -164
rect 1064 -198 1160 -164
<< nsubdiffcont >>
rect -1064 -198 1064 -164
<< poly >>
rect -1000 95 1000 111
rect -1000 61 -984 95
rect 984 61 1000 95
rect -1000 14 1000 61
rect -1000 -112 1000 -86
<< polycont >>
rect -984 61 984 95
<< locali >>
rect -1160 164 1160 198
rect -1160 -164 -1126 164
rect -1000 61 -984 95
rect 984 61 1000 95
rect -1046 2 -1012 18
rect -1046 -90 -1012 -74
rect 1012 2 1046 18
rect 1012 -90 1046 -74
rect 1126 -164 1160 164
rect -1160 -198 -1064 -164
rect 1064 -198 1160 -164
<< properties >>
string FIXED_BBOX -1143 -181 1143 181
<< end >>
