magic
tech sky130A
magscale 1 2
timestamp 1698067942
<< pwell >>
rect -1196 -229 1196 229
<< nmos >>
rect -1000 -81 1000 19
<< ndiff >>
rect -1058 7 -1000 19
rect -1058 -69 -1046 7
rect -1012 -69 -1000 7
rect -1058 -81 -1000 -69
rect 1000 7 1058 19
rect 1000 -69 1012 7
rect 1046 -69 1058 7
rect 1000 -81 1058 -69
<< ndiffc >>
rect -1046 -69 -1012 7
rect 1012 -69 1046 7
<< psubdiff >>
rect -1160 159 1160 193
rect -1160 -159 -1126 159
rect 1126 -159 1160 159
rect -1160 -193 -1064 -159
rect 1064 -193 1160 -159
<< psubdiffcont >>
rect -1064 -193 1064 -159
<< poly >>
rect -1000 91 1000 107
rect -1000 57 -984 91
rect 984 57 1000 91
rect -1000 19 1000 57
rect -1000 -107 1000 -81
<< polycont >>
rect -984 57 984 91
<< locali >>
rect -1160 159 1160 193
rect -1160 -159 -1126 159
rect -1000 57 -984 91
rect 984 57 1000 91
rect -1046 7 -1012 23
rect -1046 -85 -1012 -69
rect 1012 7 1046 23
rect 1012 -85 1046 -69
rect 1126 -159 1160 159
rect -1160 -193 -1064 -159
rect 1064 -193 1160 -159
<< properties >>
string FIXED_BBOX -1143 -176 1143 176
<< end >>
