** sch_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/tt05_analog_test.sch
.subckt tt05_analog_test VPWR VGND ua[0] ena clk rst_n ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
*.ipin VPWR
*.ipin VGND
*.iopin ua[0]
*.ipin ena
*.ipin clk
*.ipin rst_n
*.iopin ua[1]
*.iopin ua[2]
*.iopin ua[3]
*.iopin ua[4]
*.iopin ua[5]
*.iopin ua[6]
*.iopin ua[7]
*.opin uo_out[0]
*.opin uo_out[1]
*.opin uo_out[2]
*.opin uo_out[3]
*.opin uo_out[4]
*.opin uo_out[5]
*.opin uo_out[6]
*.opin uo_out[7]
*.ipin ui_in[0]
*.ipin ui_in[1]
*.ipin ui_in[2]
*.ipin ui_in[3]
*.ipin ui_in[4]
*.ipin ui_in[5]
*.ipin ui_in[6]
*.ipin ui_in[7]
*.ipin uio_in[0]
*.ipin uio_in[1]
*.ipin uio_in[2]
*.ipin uio_in[3]
*.ipin uio_in[4]
*.ipin uio_in[5]
*.ipin uio_in[6]
*.ipin uio_in[7]
*.opin uio_out[0]
*.opin uio_out[1]
*.opin uio_out[2]
*.opin uio_out[3]
*.opin uio_out[4]
*.opin uio_out[5]
*.opin uio_out[6]
*.opin uio_out[7]
*.opin uio_oe[0]
*.opin uio_oe[1]
*.opin uio_oe[2]
*.opin uio_oe[3]
*.opin uio_oe[4]
*.opin uio_oe[5]
*.opin uio_oe[6]
*.opin uio_oe[7]
* noconn ua[2]
* noconn ua[3]
* noconn ua[4]
* noconn ua[5]
* noconn ua[6]
* noconn ua[7]
* noconn rst_n
* noconn clk
* noconn uio_in[0]
* noconn uio_in[1]
* noconn uio_in[2]
* noconn uio_in[3]
* noconn uio_in[4]
* noconn uio_in[5]
* noconn uio_in[6]
* noconn uio_in[7]
xdac VPWR dac_int ui_in[2] ui_in[1] ui_in[0] VGND dac
xringosc VPWR ro_int ui_in[6] VGND ringosc
XR1 uio_oe[0] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR2 uio_oe[1] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR3 uio_oe[2] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR4 uio_oe[3] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR5 uio_oe[4] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR6 uio_oe[5] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR7 uio_oe[6] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR8 uio_oe[7] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR9 uio_out[0] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR10 uio_out[1] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR11 uio_out[2] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR12 uio_out[3] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR13 uio_out[4] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR14 uio_out[5] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR15 uio_out[6] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR16 uio_out[7] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR18 uo_out[1] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR19 uo_out[2] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR20 uo_out[3] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR21 uo_out[4] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR22 uo_out[5] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR23 uo_out[6] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR24 uo_out[7] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR17 uo_out[0] VGND VGND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
* noconn ena
xtgro VPWR ua[0] ro_int ui_in[5] VGND tg
xtgdac VPWR ua[1] dac_int ui_in[3] VGND tg
xtgbyp VPWR ua[0] ua[1] ui_in[7] VGND tg
* noconn ui_in[4]
.ends

* expanding   symbol:  dac.sym # of pins=6
** sym_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/dac.sym
** sch_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/dac.sch
.subckt dac vdd vout in2 in1 in0 vss
*.ipin vdd
*.ipin vss
*.opin vout
*.ipin in0
*.ipin in1
*.ipin in2
xdrv_b2 vdd in2 v2 vss dac_drv
xdrv_b1 vdd in1 v1 vss dac_drv
xdrv_b0 vdd in0 v0 vss dac_drv
XR1 net6 vout vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
xdrv_dummy vdd vss net4 vss dac_drv
XR2 net1 v2 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR3 vout net1 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
.save v(vout)
.save v(v2)
.save v(v1)
.save v(v0)
XR4 net5 net6 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR5 net7 v1 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR6 net6 net7 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR8 net2 v0 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR9 net5 net2 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR10 net3 net4 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR11 net5 net3 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XRDummy1 vss vss vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XRDummy2 vss vss vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
.ends


* expanding   symbol:  ringosc.sym # of pins=4
** sym_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/ringosc.sym
** sch_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/ringosc.sch
.subckt ringosc vdd clk_out ena vss
*.ipin vdd
*.ipin vss
*.opin clk_out
*.ipin ena
.save v(ph1)
.save v(ph2)
.save v(ph3)
xro1 vdd ena ph1 ph2 vss ringosc_delay
xro2 vdd vdd ph2 ph3 vss ringosc_delay
xro3 vdd vdd ph3 ph1 vss ringosc_delay
xbuf1 vdd ph1 net1 vss ringosc_buf
xbuf2 vdd ph2 net2 vss ringosc_buf
xbuf3 vdd ph3 clk_out vss ringosc_buf
* noconn #net1
* noconn #net2
.save v(ena)
.ends


* expanding   symbol:  tg.sym # of pins=5
** sym_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/tg.sym
** sch_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/tg.sch
.subckt tg vdd s1 s2 tgon vss
*.ipin vdd
*.ipin vss
*.ipin tgon
*.iopin s2
*.iopin s1
XM3 s1 tgon s2 vss sky130_fd_pr__nfet_01v8 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4A s1 tgon_n s2 vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4B s1 tgon_n s2 vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 tgon_n tgon vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 tgon_n tgon vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  dac_drv.sym # of pins=4
** sym_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/dac_drv.sym
** sch_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/dac_drv.sch
.subckt dac_drv vdd in out vss
*.ipin vdd
*.ipin vss
*.ipin in
*.opin out
XM1 net1 in vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2A net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4A out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out net1 vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2B net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4B out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ringosc_delay.sym # of pins=5
** sym_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/ringosc_delay.sym
** sch_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/ringosc_delay.sch
.subckt ringosc_delay vdd ena in out vss
*.ipin vdd
*.ipin vss
*.ipin in
*.opin out
*.ipin ena
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 L=10 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2A out in net1 vss sky130_fd_pr__nfet_01v8 L=10 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMcap1 vss out vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMcap2 vdd out vdd vdd sky130_fd_pr__pfet_01v8 L=2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2B net1 in vss vss sky130_fd_pr__nfet_01v8 L=10 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMpowerdn in ena vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ringosc_buf.sym # of pins=4
** sym_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/ringosc_buf.sym
** sch_path: /home/jakob/Documents/tt05-analog-test-main_v4/xschem/ringosc_buf.sch
.subckt ringosc_buf vdd in out vss
*.ipin vdd
*.ipin vss
*.ipin in
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2A out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2B out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
