magic
tech sky130A
magscale 1 2
timestamp 1698067942
<< nwell >>
rect -296 -1184 296 1184
<< pmos >>
rect -100 -1036 100 964
<< pdiff >>
rect -158 952 -100 964
rect -158 -1024 -146 952
rect -112 -1024 -100 952
rect -158 -1036 -100 -1024
rect 100 952 158 964
rect 100 -1024 112 952
rect 146 -1024 158 952
rect 100 -1036 158 -1024
<< pdiffc >>
rect -146 -1024 -112 952
rect 112 -1024 146 952
<< nsubdiff >>
rect -260 1114 260 1148
rect -260 -1114 -226 1114
rect 226 -1114 260 1114
rect -260 -1148 -164 -1114
rect 164 -1148 260 -1114
<< nsubdiffcont >>
rect -164 -1148 164 -1114
<< poly >>
rect -100 1045 100 1061
rect -100 1011 -84 1045
rect 84 1011 100 1045
rect -100 964 100 1011
rect -100 -1062 100 -1036
<< polycont >>
rect -84 1011 84 1045
<< locali >>
rect -260 1114 260 1148
rect -260 -1114 -226 1114
rect -100 1011 -84 1045
rect 84 1011 100 1045
rect -146 952 -112 968
rect -146 -1040 -112 -1024
rect 112 952 146 968
rect 112 -1040 146 -1024
rect 226 -1114 260 1114
rect -260 -1148 -164 -1114
rect 164 -1148 260 -1114
<< properties >>
string FIXED_BBOX -243 -1131 243 1131
<< end >>
