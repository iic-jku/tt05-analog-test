magic
tech sky130A
magscale 1 2
timestamp 1698067942
<< nwell >>
rect -246 -1184 246 1184
<< pmos >>
rect -50 -1036 50 964
<< pdiff >>
rect -108 952 -50 964
rect -108 -1024 -96 952
rect -62 -1024 -50 952
rect -108 -1036 -50 -1024
rect 50 952 108 964
rect 50 -1024 62 952
rect 96 -1024 108 952
rect 50 -1036 108 -1024
<< pdiffc >>
rect -96 -1024 -62 952
rect 62 -1024 96 952
<< nsubdiff >>
rect -210 1114 210 1148
rect -210 -1114 -176 1114
rect 176 -1114 210 1114
rect -210 -1148 -114 -1114
rect 114 -1148 210 -1114
<< nsubdiffcont >>
rect -114 -1148 114 -1114
<< poly >>
rect -50 1045 50 1061
rect -50 1011 -34 1045
rect 34 1011 50 1045
rect -50 964 50 1011
rect -50 -1062 50 -1036
<< polycont >>
rect -34 1011 34 1045
<< locali >>
rect -210 1114 210 1148
rect -210 -1114 -176 1114
rect -50 1011 -34 1045
rect 34 1011 50 1045
rect -96 952 -62 968
rect -96 -1040 -62 -1024
rect 62 952 96 968
rect 62 -1040 96 -1024
rect 176 -1114 210 1114
rect -210 -1148 -114 -1114
rect 114 -1148 210 -1114
<< properties >>
string FIXED_BBOX -193 -1131 193 1131
<< end >>
